O      �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �I]    �I]    �j& �	                   �	                      OS.iso                                                                                                                                              8�և�                                                                         �.G             6+Շ�  �%�A                          ��p     �$r                                                   �$r             �       ��b��                         �p                        ����        y��vj-  ~�b��   �p             Yj��          ���vj-  ~�b��  `J             Yj��  8                              �b��                          Yj��  ��vj-  ~�b��  ��p             Yj��  8                              �b��                                 !"#$%&'()*+,-./                                      �me��     �  0�i��         xyz{|}~0�i��  d�e��  
       0�i��  ��p     
       �����������������     �me��  0�i��  ��p     �XJ     ��������0�i��  �ne��          �XJ            MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  d� E�	] � .x  � '   
  �    �       @                         `    g�&                                                 � �           0 ��                                          @{
 (                   �� p                          .text   ��	      
                ` P`.data   �.   
  0   
             @ `�.rdata   �   @
  �   6
             @ `@.pdata  ��   0  �                @ 0@.xdata  t�   �  �   �             @ 0@.bss    @   �                     � `�.idata  �   �     �             @ 0�.CRT    p         �             @ @�.tls              �             @ @�/4         0     �             @ PB/19     F�  @  �  �             @ B/31     �   �     \             @ B/45     m   �     v             @ B/57     `        �             @ @B/70     �         �             @ B/81     �   0     �                    @ B/92     �   P     �             @ B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �D  f.�     H��(H�u�
 1��    H�v�
 �    H�y�
 �    H�<�
 �    H��
 f�8MZtXH��
 ��� � ��t5�   ��^ �V_ H���
 �����  H�Ox
 �8tZ1�H��(� �   �^ ��@ HcH<Hȁ8PE  u��Hf��t9f��u����   �z������   1҅����h���H���  脠  1�H��(Ãxt�K���D���   1�E�����7���D  f.�     H��8H�%�
 L�ξ H�Ͼ H�о � ��� H��� H�D$ H���
 D���] �H��8��    AUATUWVSH��   1��   H�T$ H���H�H�=ȃ
 D�E����  eH�%0   H�܂
 1�H�pL�%+� �H9��4  ��  A��H���H�3H��u       �H�5��
 1����"  ����q  ��    ����  ���1  H��
 H� H��tE1��   1����D�  H���  ��� H�0�
 H�舦  H������<] ��  H���
 H��� �4] 1�H� H��u�_�     ��t,��t'�   H����� ~�A��A����"AD���fD  ��u�f.�     �� H�����u�H�1� D�E��t�D$\�
   ��   ���	 �� D�cMc�I��L����Z ��H�=� H��~K�C�1�L�,�   �    H��GZ H�pH����Z I��H�D H�H��H���Z I9�u�J�D%�H�     H�-�� 趚  H���
 H�h� �r� H� H�L�U� H�V� �  �;� �9� ����   �#� ��u�N[ �� H�Ę   [^_]A\A]��D$`����fD  H�5��
 �   ���������   �[ ��������H���
 H���
 �Z ���   �����1�H������f�     H����� �6���f�H���
 �   H�l�
 �gZ �{������Z �f.�     H��(H���
 �    �ʙ  ������H��(�@ f.�     H��(H���
 �     蚙  ������H��(�@ f.�     H��(��Y H��������H��(Ð������H�	   �����@ Ð��������������UH��H�� ��  H��*
 H�%y
 ��	 H�)y
 H���!Z ��X �    H�� ]�UH��H�� H��� �MR	 �H�� ]�UH��H�� �M�U�}u!�}��  uH�b� �]J	 H������1����H�� ]�UH       ��H�� ���  �   �����H�� ]Ð�����������UH��H�� H�!� ��Q	 �H�� ]�UH��H�� �M�U�}u!�}��  uH�� ��I	 H����������H�� ]�UH��H�� ���  �   �����H�� ]Ð�����������%�� ���%^� ���%N� ���%n� ����OweL��F
 ��Ic�L���f�     M��tED�Q(D;Q,};Ic�A��L�@H�A J���@    D�Q(�L�@L�H��     M��tM��u�1�� L�IE�I��A��RtA��Ot	H���D  D�YHA��R�    A�Cu	A�C�   I���AHL�IE1��A����UWVSH��(M��H��H��L��t#H�5G
  �;Ow�Hc�H���H�[H��u�H��([^_]�H�[���     L�CA�8u�E L�CH��H������H�[���L�C��@ UWVSH��(M��H��tpH��   J�,H���"H��H��H��H��   H9�@�<@��  t>H=�   �>uӺ�   ƃ�    L��  H����  �   1҃�@  ��    H��([^_]��    VSL�	E�A��n�}   A�@�<	��   1�I��E1Ҿ���A������A�@Љ�I��)�A����D9�|2C��L�	A�@E�D�P�A�PЀ�	v˺0   )�DE�D��[^� A�����D��[^�@ I�AH�E�AA�PЀ�	wI���   �o���E1���f�     SH�� �A(;A,}7HcЃ�H��L�RH�QJ���C    �A�A   �����CH��H�� [�1�H��H�� [ÐSH�� H�Q�H��<_t-<nt-H�I�������xH�S�:_uH��H�SH�� [�@ 1���������D         SH�� H�A�8TH��uOH��H�A��������x<�S(;S,}4Hc�L�@H�C J���@    �S(�    �HH�� [�f�     1�H�� [��     SH�� H��H�I����1҅�~sL�KHc�H�KL)�H9���   L��CH�St	�:$��   ��	�K(�S,D9���   Hcу�M��L�RH�S J���B    �K(txH�    L�J�BH�S@H��H�� [�I�_GLOBAL_M9u&E�YE�C�A��;wI�     M��sA�y	NtH9�}$Hcу�L�RH�S J���B    �K(�fD  1��H����	�K(H�S�S,�D���� D�SHE�BA)�9�D�CH}�Hc���H�@H�C �K(H��H�QD
 H�    H�B�B   �0���f.�     WVSH�� H�AH�y@�8BH��H��u5fD  H��H��H�C�p���I��K   H��I������H��H�C�8Bt�H��H�{@H�� [^_�f�VSH��(H�A�8SH��ucH�HH�K�x u`1��KE1Ƀ�A��u��tH�S���C���   DFʹt   H��O
 L���  ��
8���   H��8L9�u�1�H��([^�f�H�HH�K�@�HЀ�	w1�<_u&9K8v�H�C0H��H��([^�f�<_t��H����b����H�1Ҁ�	w3fD  �ҍL��9�w�H�C�8 t<H�PH�S� <_t�ʍHЀ�	vӍH����l����ҍL���Ń��f�     1�����f.�     L�R(�K(D�C,M��t;D9�D�Z0��   Hc���H�4@H�C H���@    �K(�    L�PD�XH�C@E��t{L�J�R SHD9�}uHc���L�@H�C J���@    �K(�    L�H�PH�S�:B�����H��       H�������H��������S8;S<�����H�K0Lc�J���S8�|���L�J�R�1��1��h����VSH��(��H��uH�A�8 u
1�H��([^ÐH�PH�Q���htD��vu�H�sH������H�C�8_u�H��H�C�	���H�C�8_u�H��H�C�   H��([^�H�K������ؐ��P���'v<Dt1��H�  �   ��H�����Q�B�<����߀�O��	����SH�� H�A�8_H��uH�PH�Q�x_t!H�I�x�����1���x�   H�� [�D  H�IH��H��P�����x��	~�H�S1��:_u�H��H�S��1���@ f.�     H��t �9/u����9/u��tH�I��H��u�1��u�H�AÐH��   H��t�H�@��H�Hx�@ ǁ0     1�H���WVSH�� H��H��H��t>H�5@
 �;Kw�Hc�H����    H�SH�������H��uH�[H��u�fD  1�H�� [^_�fD  H�SH���d���H��t߃8/u�H�� [^_�f�UWVSH��(I�@I�pH�DH��H��A�PH9�L��w9��u#H�KI��H��H�M H�H�HC�  H{H��([^_]�f�     ��u�H��t+�    H�H9�w�H�H���%M H��tH��SH�s�H���   w���H��M H�    H�C    H�C    �C   ��    SH�� H�A�8LH���  H�PH�Q�H��_�  ��Z��   H���u  H����   �8'�  L�S�<   A�
��nuI�RH�SA�JI�Һ=   ��E�  ����   I�J�D  H��E����   H�KD�	A��Eu�D)�D�C(D;C,��   Mc�A	       ��M��O�IL�K O��A�A    D�C(��   ����   I�    M�QA�IH��I������H�S�
��EuH��H�SH�� [�1�H�� [��     ��_tH��H��H�S1��"  H�S�
�H�PH�S�H��Zt�1��H�P�J��������R)SH������E1��s���1������AUATUWVSH��(H�Q�H��<L��  <T��  <s��   <ft>�HЀ�	�s  H���  H��H���3  H�C�8I��  H��H��([^_]A\A]Ð�zptzH����  H��H����   � ��1�L  ��2��  ��3��   H�C�8_�r  E1��:  @ �B<r�d  <pu�H��H�Q�#���E1ɺJ   I���.   H�BH�A�zT�~  �����������������tk�S(;S,}cHcʃ�L�IH�K J�4��F    �S(�   �F����<it<t�����zl����1�<t��  H���  H�SH�ƀz ��  1�H��H��([^_]A\A]�f�     H��([^_]A\A]����<ou��zn�����H��H�S�r���@ H��([^_]A\A]�_���H�UH�=�<
 �   �BL�"��CHL����� ���q  D�jA����  �M  A����  A���N���H�=Y<
 �   L����� ���P  A�$<f��  <n����A�D$<wt<a�	����_   H���  H��H���  H��H�C���E��  ��p��  ��i������xl�����H���5���I��I���;   H���2���I��:   I���"���I��9   I��� D  H��H��H�C�@  I��   I��H��H��([^_]A\
       A]������H��H�Q��
  H��H���  H��H�C�8It/I��I��   �H��H��H�S�E   �*  I��0   I���H��H��H�C�  I���   H��I���j���I��   I���e���f.�     A�$<p��   <m��   E1�H�=�:
 �   L����� ����   H������E��tI��I���8   H�������I��I��6   �����H���E   H��H�C�e  �� �E���L  �3������+���E1�I��5   ����fD  E��t�1�����@ H��1�H�Q�����A:D$�:���H�C�8_�0���H��H�C� ���H���  �<���H�EH� �xc�  A�<$f�3  H������I��H�=�9
 �   L����� ����   H�=�9
 �   L����� ��tH�=l9
 �   L����� ����   H���  H��H�C�8I��   I��M��8   H������I��7   I������fD  H���  I��6   I������H���`����q���H���S���H��H���H���H��H���=���H��I�������1������ �P���v��r<�����H���,  I��������E   H���   H���F���H���7  I�������H�������H���&���H���  �o���H��H��H�C�  I��   H��I������H��������xi����H���E   H��H�C�   I���>���H��E1�H�C�.���UWVSH��8H�A8H�t$(H�ˉ�H�D$(    u'�kE1ɺ.   H���;���H��H�t*H�pH�C@8(t(�{LH���CL   ����H��I���{Lu�1�H��8[^_]�H��H�CH�D$(H       ��8[^_]��     H��E1�E1��.   H�AH��8[^_]�����UWVSH��8H�QH�q@�H��<E��   H�D$(    H�|$(�Hf���I<��   H����   I��M����   E1ɺ/   H���a���H��H�tiH�SH�x�<Etj<Lt9~�<Xu@H���kLH���CL   H�S����I��H�C�kL�8Eu'H��H�C�H���e���I���H���  I���v���1�H��8[^_]�D  H�D$(H��H�s@H�SH��8[^_]�fD  H��E1�E1�H�Q�/   H��8[^_]����H�Q���I<wH��H�Q�����D  1�� f.�     AUATUWVSH��HH�Q�H��<S��  ��   <U�	  <Z��  H��H�Q1��}  H��H���X  H�C�8E�K  H�PH�S�P��s�  ��d�F  H���~���H��I��t� �����E��  �>��  I��   H������H����   �    <N�  H��A�   H�QH�T$8�P  H��H����   1�H��E1������H�SH��    I���2@����   @��D�   �N�H��H�����&�    C��N����~  ���v  @��S��  @��I��  @��T��  @��E��  M��t(@��Mu"H�BH�C�JH�� ���v���f�     H�    1�H��H��H[^_]A\A]��    �zt��   1������H��H�C�8Iu��3�H���h  H��H�C�8Iu�H��t��C8;C<}�H�S0Hcȃ�H�4ʉC8H������I��   H��I���C���H���t����  H��H��H��H[^_]A\A]� H��H�Q��  �S(;S,I����  H�C Hcʃ�H�       I�S(L��H��3
 I�     I�@A�@   �   H��������CHH��H�C�8I������3���H���  M����   I��H�S@��S�
�������E��   M��������C8;C<�����H�K0Lc���N�,��C8�
���������BH�ك��<T�~   �I  M��   u/H�SI���
� M���G���H��H��H�S�G����   f�M��I��H�������I���O���f.�     �   ��f�     �E   �v���fD  �  �}���fD  H��H��H�C�������������H������H��H��t� �����E�d  �C(;C,�C  HcЃ�H�RH�S L��A�A    �C(A�F   A�iI�y�c���M��L�/�f���M��tH�D$8L�d$8I�D$�:E�I���H��H�t$8H�S�9���H�F�8)�$���H�@    ����fD  H��H��H�C� �����������C(;C,��   HcЃ�H�RH�S �C(H�.1
 L��I�    I�AA�A   �����     �   H�������M�������H�SI���
�������f�     E1��s���H��L�L$(�k���L�L$(���e����Q���E1��I���H���I��������H���<�����������6���D  f.�     ATUWVSH��0L�AH��L����������   A��A�<JwdH�q0
 ��Hc�H����sLH���CL   ����E1ɺB   H��I���sL����H��H�D$(tH�S�: tH�JH�K�:E��   D  1�H��0[^_]A\� H�T$(E1�H���   H��H��t�H�CH�ـ8Ft`�7���H��H�H��t��:H�D$(�O��wH�JH�BH�H�       D$(H�H�D$(H��t��S8;S<}�H�K0Lc�J���S8H��0[^_]A\��7  H��H��H���G���H�D$(f�H���G����S8;S<�;���H�K0Lc�J��H�D$(�S8H��0[^_]A\�f.�     I��H��L�C� ���E1ɺ(   H��I���M���H�D$(�fD  H�iD
 �ыK(��aHc�H��H�;K,�p�	 Hc�I����L�@H�C J���@    �K(H�P�R� '   SHL�C����@ I��H��L�C�p���H�D$(H��H�C�8I��  H�������I��!   H��I������H�D$(�����fD  H������H�sH�D$(�>I������SP���  H�������S8;S<�����H�K0Lc�E1�J���S8��P���wH��H�sH���g���I��L�D$(�   H������H�D$(�X����     A�@��0</�   H������  H����  1�H���2���H�SH�D$(�:I�b���H��H�S�fD  I��H��L�C����E1ɺ#   H��I������H�D$(����� I��H��L�C����E1ɺ&   H��I���]���H�D$(���� H���  H�D$(����I�@H�CA�x �����I�@H�CA�@��F<0�����H��-
 ��Hc�H���I��H��L�C� ���E1ɺ%   H��I�������H�D$(�#��� I��H��L�C�����E1ɺ"   H��I������H�D$(����� I��H��L�C����E1ɺ$   H��I���}���H�D$(����� M�HL�KA�@<_��  ��0L��<	v�  H��H�QH�S�A��0<	v�I�ҋC(M)�;C,�����Lc���E��O�@L�C K�4��F           �C(�����H�    L�ND�V�A<_I��������I��H��L�K�����I��*   H��I������H�D$(���� I��H��L�C����H��H���4���H������H��I��� ���I��+   H���p���H�D$(����A�x_�u  H�������H��H�������H�C�8_�����H��H��H�C�:���I��-   H��I������H�D$(�]����S(;S,���	 H�=�C
 Hc�H�@H�C H���@    �S(� '   H�x�CH�m����S(;S,���	 H�=�C
 Hc�H�@H�C H���@    �S(� '   H�x�CH�+����S(;S,�<�	 H�=�C
 Hc�H�@H�C H���@    �S(� '   H�x�CH������S(;S,�����H�=�)
 Hc�H�@H�C �S(H��H�     H�x�@   ����H������E1ɺJ   H��I�������H�D$(�3����S(;S,�J�	 H�=�B
 Hc�H�@H�C H���@    �S(� '   H�x�CH�C����S(;S,�A�	 H�=>B
 Hc�H�@H�C H���@    �S(� '   H�x�CH
�����S(;S,���	 H�=�A
 Hc�H�@H�C H���@    �S(� '   H�x�CH	�����S(;S,���	 H�=�A
 Hc�H�@H�C H���@    �S(� '   H�x�CH	�}����S(;S,�o���H�=e(
 Hc�H�@H�C �S(H��H�     H�x�@   �>����C(;C,���	 HcЃ�H�RH�S H�4�1��F    �C(H�t$(�,   A�@��0<	��f�VwH�K����H�t$(H���N���H�FH�D$(H�x �����H�K�����H�C1Ҁ8 tH�PH�       S�H�D$(��s����f�P����@ H���x���H��H�D$(�z����8�*����n���1������H��H��H�C�����L�D$(�   H��I������H��H�D$(������{LH���CL   �q���H��H�Ɖ{L����H�S��z���H�FH��D�c(H�C�k8�{H����H�S�:ItH�sH�D$(D�c(�k8�{H�{���L�D$(M��������S8;S<�����H�K0Lcʃ�N��I��H�ىS8�   �����H�D$(�6����{LI��H���CL   L�C����H�Ɖ{L�q����VSH��(H�A�8 H����   H�PH�Q�x D���   1�L�4
 A�C   1� D��)щ�������Hc�H�IM��I�	D8t~[A��D9�u�1�H��([^�f.�     @8qu݋S(;S,}�Hc�H�@H�C H���@    �S(� 1   L�HH��([^�D  �P�E1��_��� H�PA��vH�Q�pu^�F�<	�A����n����S(;S,I���l���H�C Hcʃ�M��H�IH���@    �S(�G���@��H� 2   ��0L�@�P�/���A��c�����@��v������QL1��qP�����AP�g����KPE1�I����t�4   H���=����sPH��([^ú3   H���&�����@ VSH��8H�QH�D$(    �H��<EA������A�ulH�t$(<.����t@�\�    E1ɺ.   H�������H��H�t=H�SH�p���A��<E��A�u-<.t)<Rt<Ou�zEtH������H��I��u�1�H��8[^�f�H�D$(H��t�H�x u�H�P�:'u�H�R�z	uӋR)SHH�@    ��f�f.�     AWAVAUATUWVSH��(E��L�AH��H��A��H��E�A       ���A��A��L��E�E�A���A��A�����������������   f�I�@A��rH�C��   A��V�  A��K�  A�x tfI�@H�CA�@<x�  ��߀�O�  �CH	<O�D  D�{LH���CL   �a���H��I��D�{LtH�C�8EuH���N   H�C�&1�H��H��([^_]A\A]A^A_��    �CH	��E1�E1�H������H��H�t�L�CH�pL��E������������A��u�A��Ft�f.�     ����   H��H9�t�H�?�����   ��u��   �� �CH	D��E1��z�����CHD��E1��j�����CHE1ɺL   �X���<w�*����CHH���K���H��I������H�C�8E����H���O   H�C����E1ɺN   ���� �   �N���D  �   �>���D  VSH��(H�A�8JH��t^��t:H������H��H��t<H�������H��I��t,I��)   H��H��([^�����@ H��1�����H��I��u�1�H��([^�D  H��H�A�fD  SH�� H�A�8FH��uOH�PH�Q�xYt1�   H���T���H��H�������H�S�:Eu H��H�SH�� [�f�H��H�A��fD  1�H�� [��     UWVSH��(H��H�I��PЀ�	��   �P���w<<o��  H���*���H��H��t	�81��   H�C� <B��   H��H��([^_]ÍP�����  <L�  <U�<  �A<l��  <t�(  H�A1�H�C�A<tu�H��H�KH���L�����x��S(;S,�=  Hcʃ�L�IH�K J�,��E    �S(H�S�E�C8;C<�E G   �N  H�K0Lc       ���J�,��C8��;���H������H��H�C� <B�)���H��H��H��([^_]�����H�@H�=y!
 �KH�PH�0�T�   �SH��� �������H���I���I��6   H��I������H������H��H�KH������H��H��tH�������������1�H��H��([^_]��     �yn�T���H��H�K�G���f�     H�S@H��tD�E����   A����   <D��   �A<I��  ��1<w�L��'
 ��H��A�4�H�K�C(;C,��  Hcȃ�H��L�IH�K J�,��E    �C(��  �F�����  H�E    �uH�U�����BCH�<C�u���<D��   �A��0<����L� 
 ��Ic�L���A�   H�AH�C�C(;C,}^Lc���H��O�@L�C K�,��E    �C(t=H�E    D�UH�U�A�2���A�   �A�   �A�   �A�   �@ �A1�����D  H�A1�H�C�A<l�����H��H�KH������H��H�������H�S�<E�����H��H��H�S�_�����x\�S(;S,L�C��   Hcʃ�L�IH�K J�,��E    �S(�E�C8;C<�E E   H�u}kH�S0Hcȃ�H�,ʉC8A� �M���H�C1�� �?���H�AH�C�A��1<w;H��%
 H����H�KH�ً4������H�S@������1������A� 1�������A1�������     WVSH�� H�A���H�ˀ�Gtx��Tts����H��H���d  ����   �C��   � �P��3�R  H�      H��s&A�   H��H�v��H��3�'  L��H��H��u�H��H       �� [^_Ð�KH�Q�SH���T��  ��G��   H�PH�S�x ��   H�PH�S�x�W���1��   H��
 ��Hc�H���D  H�C� ��t�<Et�H���� ��   ����   ����  ����   H�BH��tS���4wLI��     �   H��L����   ��A�   u�$���4wL��H��L����   ��t	H�@H��uܺ   �   H�s1�H��H�� [^_Ð�������H�V�����3�����H�      H�������A�   H��H�R�:�O��3wL��H��H��u�H�V����fD  ��Lt
r��N��wH�RH�������@ 1�H���v���H��I���\�����u�>u�8)uH�@    @ I��   H��H�� [^_�I���f�     H�PH�S�x ����H�PH�S�@��C<3�����H��
 ��Hc�H���@ H������E1ɺ   I��듀x tH�PH�S�xn��  1�H������E1ɺH   I���a���f�     H���8���H��H���-���I��   I���5���1�H�������E1ɺ   I������ H�K�7������@���H�S�: �3���H�rH�s�:_�"����x�E1����������$��  �F<S�  <_�  <$������$   H�s�C(H��;C,�����HcЃ���L�RH�S N��A�A    �C(A�@   A�IH�sM����  �?   H������H��I����������^���E1ɺ>   �3���H������E1ɺ   I������ H�������E1ɺ   I��� ����     H���X���E1ɺ   I��������            H���8���H�KH��������������H�C�8_�����H��H��H�C����I��   �CHI������ �v   H���C����������1�H������E1ɺ   I���Y�����h   H���������}���1�H�������E1ɺ   I���)����1�H����������P���1�H����������>���1�H������E1ɺ   I�������f�H�������E1ɺ   I��������     ���KHH���"���E1ɺ	   I������f���
�KHH������E1ɺ
   I������f�H�������E1ɺ   I���p����     H�������E1ɺ   I���P����     H�R������    �   �f�     �L�J��$t��t
L��9�A���C(;C,}gHcȃ�D)�L�IH�K N��A�A    �C(I�    I�qH�sE�QH�H�s�\���M���v���fD  �.   ����fD  �/   �����HS1�����1�H���1���E1ɺI   I���y����AWAVAUATUWVSH���   M��H��A��L���[  D��0  E���  A���O�O  L�L
 ��Ic�L���H�E�88�   L�EI�@H� �xc��6  L�MD��H����V  ����  H�E�81��=  H�@L�%�
 �   L��H�UH�0L�B��� ��u
A�8��?  D��H���U  L�EH�=
 �   I�@H�H����� ���]:  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H��H�PH��   D���[ƃ  [H�EL�@��@  H��   �   u.ƃ�    L��  ��   H����  Hǃ              ��@  H��   H�PH��   �]ƃ  ]H�E�81ukH�@�xuaH�@�8>uXH��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �)ƃ  )H���   [^_]A\A]A^A_�I�QH��A�   L��   H��   H�P�A���H����6  L��   �ǃ0     �@ ǃ0     �H�UH��E1��5���H��u�w;  A�ԃ8/�8&  H�x �-&  H�@A�T$H��u�L�}D�d$(A��H�-�
 ��A��E9��:���D��<  M��D��H���?  D;t$(}�H��   H�=�
 �,   �'f�H��H��H��H��   H9�@�4@��  t��7H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  �H�5	
 H��   �n   L�f�)H��H��I9�H��   @�<@��  ��"  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5v
 H��   �{   L�f�1�     H��H��I9�H��   @�<@��  �!  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �{   L�f�3f.�     H��H��H��H��   I9�@�<@��  �F"  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5O
 H��   �g   L�f�3f.�     H��H��I9�H��   @�<@��  ��!  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �g          L�f�3f.�     H��H��I9�H��   @�<@��  �"!  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5
 H��   �d   L�f	�3f.�     H��H��I9�H��   @�<@��  �?   �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �D�EL�d$@H��
 L���S L��
H����������!�%����t�������  D�H�JHDщ� �H��L)��b���H��   I�4�&H��H��I��H��   L9�@�<@��  �/���H=�   A�<$uͺ�   ƃ�    L��  H����  �   1҃�@  �H�5:
 H��   �t   L�f�/fD  H��H��I9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H��   �uH�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   @�4@��  �#���L�ED��H���:  L�ED��H����9  � ���H�5�
 H��   �j   L�f�)H��H��L9�H��   @�<@��  �#  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H�ٿ    H�5�
 L�f�d9  H��   �)H��H��H��H��   I9�@�<@��  �  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�E1��8'�%  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H��H�       PH��   D���(ƃ  (L�E�8  H��   H=�   �q)  H�PH��   �)ƃ  )�} =��*  ����)  L�ED��H���=8  �?���H�E�8:�{���H�@�8;�n���L�EL�MD��H���KM  ���
���H�EH�
 L�eH�xH�@H�hH�pI�D$H�� ����5  I��D��H����K  M��D��H���3K  I��D��H����K  H��A�   H�Q
 �p���I��D��H���K  ����L�eH�mA�$��1�$  ��3�F7  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H��H�PH��   D���(ƃ  (M�D$��6  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �)ƃ  )I��D��H����J  ����L�ED��H���J  ����H�5
 H��   �o   L�f�1�     H��H��L9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �o   L�f�3f.�     H��H��I9�H��   @�<@��  �7  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�mH�5
 �o   H��   L�nD�e�+f�H��H��H��H��   I9�@�<@��  ��  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �L�EH�uM��tD��H����4  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@         H��   I��D��H���{ƃ  {�4  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �}ƃ  }�A���L�EM��tD��H���&4  H�} �"���H��   H���   v+�3 H��H��1�L��  ��  Hǃ       ��@  A�,   H�=j
 L�w�*H��H��H��H��   I9�D�$D��  �2  D�'H���   u�ƃ�    ��   H�پ   L��  ��  1���@  �f�} �#  L�EH�(
 I9@��  D��H���C3  H��   H�BH���   u*��   ƃ�    L��  H����  �   1҃�@  H��   � ƃ   f�} ��  H�5j
 �_   H�n�/fD  H��H��H��H��   H9�@�<@��  ������>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H��H�l$HH��(  �D$P    H�D$@H�D$@H��(  H��   H�D$X�32  D�T$PE���B"  H�D$@H��(  ����H��(  L�d$@H�l$HH��   L��(  �D$P    H��H�L$@L��H��H�D$X�u.  H�G� �����c.  H���   ��     H�P�����w]D�pE��uL����%  L� ���H��L�D@L�@L�DHL�@L�DPL�@H�L@I�H��(  L�DX�@   H� H��u�L�ED��H���61  D�\$PH��(  E���(�����H��Iă�tM�D$��D��H��I�� �1  ��u�L��(  L�ED��H����A  �����H�5a
 H��   �n   L�f�, H��H��I       9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �h   L�f�3f.�     H��H��L9�H��   @�<@��  �  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5 
 H��   �r   L�f�3f.�     H��H��I9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5f
 H��   �T   L�f�3f.�     H��H��I9�H��   @�<@��  �Z  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �T   L�f�3f.�     H��H��L9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5;
 H��   �g   L�f�3f.�     H��H��I9�H��   @�<@��  �2  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�
 H��   �j   L�f�3f.�     H��H��I9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5
 H��   �c   L�f�3f.�     H��H��I9�H��   @�<@��  �
  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5~
 H��   �v   L�f�3f.�            H��H��I9�H��   @�<@��  �N  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  몋�8  H�E�ɋuE1����I"  ��#L��(  �,  9U �#  ��$��
  D  L�L$@H�D$@H�l$HH��(  H��   �D$P    H�D$XL�ED��H����+  �D$P���S  H�D$@E��H��(  �����L��   �����H��(  H�D$@�L��(  M��t�L���9���  H� H���g���D�@E��u�H�P�D�B�A��v�E1��F���HcUH�uH���\���H��   H�,�.�     H��H��H��H��   H9�@�<@��  �!���H=�   �>uϺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H����*  �����D�mH��   E���(  H�5�
 �{   H�n�2f�     H��H��H��H��   H9�@�<@��  ��  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �D��8  E���`  H�5L
 H��   �a   L�f�3f.�     H��H��H��H��   I9�@�<@��  �`  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �A��L��p  H��p  L��(  Hǃ(      L�EtE�E��uA�x��"  D��H���k)  ��  <�+  H��   H=�   ��  H�PH��   H��D���<ƃ  <L�E�&)  ��  >�Z  H��   H=�   �  H�PH��   �>ƃ  >L��(  L��p  �����H�EL��(  Hǃ(             H����  D�L�d$@H�D$@    H��   L��(  H�D$H�D$P    A�I��3H�T$X��  I�      I����  M�T$ A�   A�   H�@H���f  A���\  H��(  A��L��(  D�I�BA�B    I�RI�
A�I��3�i  L��I�� H��L��u�L�ED��H��H�D$(��'  H�D$(�8uH�D$0H��   D��H��L�D�^�E��u^H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  L�F�H��   H��D��� ƃ   �(  H�� I9�u�L��(  �W���L�ED��H���A'  A��H��   ��  H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �.ƃ  .H�}�?F�W  I��D��H����&  �����A��Hc}H�u��  H�������H��   H�,>�&H��H��H��H��   H9�@�<@��  �����H=�   �>uϺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H�ٿ[   H�5%�	 L�f�$&  H��   �)H��H��H��H��   I9�@�<@��  �
  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H���%  ����A��H�E�M  HchH�0H�������H��   H��&H��H��H��H��   H9�@�<@��  �a���H=�   �>uϺ�   ƃ�    L��  H����  �   1҃�@  �D��L��(  ��A�� �<  L�EM��t
A��@�4  L�E��H���.  �����H�5�	 H��   �c   L�f       �)H��H��I9�H��   @�<@��  �K  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5��	 H��   �V   L�f�0�    H��H��H��H��   L9�@�<@��  ��  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�	 H��   �v   L�f
�3f.�     H��H��L9�H��   @�<@��  �&  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H��H�PH��   D���~ƃ  ~L�E�#  ����H�5h�	 H��   �t   L�f�)H��H��I9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5�	 H��   �t   L�f�1�     H��H��I9�H��   @�<@��  ��  �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5f�	 H��   �t   L�f�3f.�     H��H��I9�H��   @�<@��  ��   �>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �L�@H�D$@L�L$@H��(  H��   H�l$H�D$P    M��H�D$X�j����a����    L�ED��H���A!  �C���L�ED��H���-!  �/���L�ED��H���!  ����L�ED��H���!  ����L�ED��H����   �����L�ED��H����   �����       L�ED��H����   �����L�ED��H���   ����L�ED��H�ٿ    H�5��	 L�f�   H��   �-�     H��H��H��H��   I9�@�<@��  t7�>H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H���   ����L�ED��H���   ����L�ED��H����  �����L�ED��H����  H��   H�PH=�   u*��   ƃ�    L��  H����  1��   ��@  H��   �]ƃ  ]����L�ED��H���y  �{���L�ED��H���e  �g���L�ED��H�ٿ-   H�5��	 L�f�A  H��   �-�     H��H��H��H��   I9�@�<@��  t7�>H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  �L�ED��H����  �����L�ED��H���  ����L�ED��H���  ����L�ED��H���  ����L�ED��H���x  �z���H�u��Q���wLH�PH=�   u.��   ƃ�    L��  H����  H�u�   1���@  H��   � ƃ   Ic�|.� uA�l$�Hc�H������H��   H��'�H��H��H��H��   H9�@�<@��  �����H=�   �>uϺ�   ƃ�    L��  H����  �   1҃�@  �H��p  H��tH��   H�D$HH�T$@H�T$@H��   L�EA�8�v  D��H���Q  H��p   �J���H�D$@H��   �9���L�ED��H���#  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��          �]ƃ  ]������EL�d$@H���	 L��D�@�l�  L��
H����������!�%����t�������  D�H�JHDщ� �H��   H��L)�taI�4�"H��H��I��H��   L9�@�<@��  t9H=�   A�<$uѺ�   ƃ�    L��  H����  �   1҃�@  �H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �}ƃ  }�����L�ED��H���  ����L�ED��H���  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �)ƃ  )�S���L�ED��H���=  �?���L�ED��H���)  �+���L�ED��H�ٿ)   ��8  H�5O�	 L�f��  H��   ��8  �%H��H��H��H��   I9�@�<@��  t7�>H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  뮋EL�d$@H���	 L��D�@�2�  L��
H����������!�%����t�������  D�H�JHDщ� �H��   H��L)�tbI�4�#�H��H��I��H��   L9�@�<@��  t9H=�   A�<$uѺ�   ƃ�    L��  H����  �   1҃�@  �H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �}ƃ  }����I��D��H���  ����L�ED��H�ً�@  �`  9�@  �[���H9�   �N���H��H��   �>���E��L�}�1���A�D$��D$(������} /L��(  �����H�������H�5��	 �_   H�n�*�H��H��H       ��H��   H9�@�<@��  ������>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�5��	 �t   H�n�*�H��H��H��H��   H9�@�<@��  �a����>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H�H9�wg����fD  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   @�,@��  H��H9������H���.H)�H��~�@��_u��~_u��~Uu�L�fL9��v���1����0��I���L9��]���A�$�HЀ�	vލH�����  ��7��HchH�pH���E���H��   H��(f�H��H��H��H��   H9�@�<@��  ����H=�   �>uϺ�   ƃ�    L��  H����  �   1҃�@  �H�UH���G���H�������8/��  H��   I��H��H�H��   D���  H��   �����EL�d$@H���	 L��D�@�'�  L��
H����������!�%����t�������  D�H�JHDщ� �H��L)��6���H��   I�4�(f�H��H��I��H��   L9�@�<@��  ����H=�   A�<$uͺ�   ƃ�    L��  H����  �   1҃�@  �L�d$@E��H���	 L���b�  L��
H����������!�%����t�������  D�H�JHDщ� �H��   H��L)�tbI�4�#�H��H��I��H��   L9�@�<@��  t9H=�   A�<$uѺ�   ƃ�    L��  H����  �   1҃�@  �H�PH=�   u*��   ƃ�           L��  H����  �   1���@  H��   �}ƃ  }����H��   ����A�   A����  H�@D�A��F�R  E�A�A��3��  H�      L���i���A��t{E��I��I��M�E�N��   L��L��(  I��A��N�T@L���K�I�J�DHH�@B�DP    J�TXD�A�I��3�  �   H��L�������I�� A��u�ǃ0     �����H�@�p����������h  �������H�E���������x�������<�����H�@� <0�G  <1�����H�N�	 A�   H���K����m���fD  H�=�	 I�D$�   �U L�0L����� ��u	���  ��8��  H�=��	 �   L���A��A�� E��E����  H�=�	 �   L����� ����
  H��M��D���W&  H�=��	 �   L����� ����  H�=��	 �   L����� �������H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   I��H��H�PH��   D���(ƃ  (�5  H��   H=�   u%ƃ�    L��  ��   H����  1���@  H�PH��   �)ƃ  )�����M�@D��H����  H��p   tH�D$@H��   H��   ��  <H����  H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   H��D���<ƃ  <H�EL�@�O  ��  >��  H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �>ƃ          >�������   ƃ�    L��  H����  �   1���@  ����H��   H���   ��  H�BH��   � ƃ   �~�����   ƃ�    L��  H����  �   1���@  ����H�5��	 H��   �_   L�f�1�     H��H��H��H��   I9�@�<@��  ������>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �I��D��H���u  ����L�E��H���r  L�EM���������H���  ����H�5��	 �:   L�f�-@ H��H��H��H��   I9�@�<@��  ������>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �H��   H���   ��
  H�BH��   � ƃ   ����ƃ�    L��  ��   H����  �)��@  ƃ  )Hǃ      �} =�m���H��   H�PH��   �-ƃ  -�K���H��   H=�   u%ƃ�    L��  ��   H����  1���@  H��H�PH��   D���[ƃ  [L�E�G  H��   H=�   u%ƃ�    L��  ��   H����  1���@  H�PH��   �]ƃ  ]�����A�������H�T$0H�T$0H��   H�D$8�����L�ED��H����  �����H���   �����ƃ�    L��  H����  Hǃ       ��@  �����H�5�	 H��   �{   L�f�%H��H��I9�H��   @�,@��  t;�.H��H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  뮋GL�d$@H��	 L��!       D�@��  L��
H����������!�%����t�������  D�H�JHDщ� �H��   H��L)�taJ�4"�"H��H��I��H��   L9�@�,@��  t9H=�   A�,$uѺ�   ƃ�    L��  H����  �   1҃�@  �H�5^�	 �}   L�f�%H��H��H��H��   I9�@�,@��  t7�.H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  �H�����A�   �����ǃ0     �����H�D$@��H��L�L$@H��(  H��   H�l$H�D$P    H�D$X�  D�|$PH�D$@E��H��(  �~���H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   � L��(  ƃ   ����I��D��H���  ����� �P���v��r<�/���D��H���_  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�ٿ>   H�5D�	 L�fH�PH��   D���<ƃ  <H�EL�@�d
  H��   �)H��H��H��H��   I9�@�<@��  ��  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  �D��X  L��P  E��~1I;�  A�J�I�QH��H���I��H��H;B���   H9�u�D;�\  ��  Ic�A��H��D��X  L�L��   H�H��M��t\Hc�h  D��l  A9���  D�AH���E�PH��E9���  E��L��`  I�qI�I�rL�M�	L��M��u�D��h  H�    H�PH��E1�蓚��H���Z����"       ��/�������<  �������H���9���H����  �����M��L��H  M�������I; t�L��H�RH�������H�
H9�t�H9�u�I9�t��x����H����W  ��W����H�ED��H��L�@�s  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �)ƃ  )������<  ���S���H���P���H���B����B���f�E1��A��H�mH��tK�} /uEH�EH��t<�8Ju�H�PH���n���1�H��u�D  H�x tH�@��H��t�8/t�A��L�d$@H���	 L���7�  L��
H����������!�%����t�������  D�H�JHDщ� �H��L)��F���H��   I�4�&H��H��I��H��   L9�@�<@��  ����H=�   A�<$uͺ�   ƃ�    L��  H����  �   1҃�@  먹   H��L����� ���P  H�ED��H��L�@��  �4���I�pH�=��	 �   ��� ������L�ED��H���s  A�   H��H���	 �>����i���L�EE�E���Z�����=��  D��H�ك��2  ���0���H���	 Hc�H���H���	 A�   H����������H���	 A�   H���ʏ�������H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �lƃ  l����H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �uƃ  u�2���H���	 A�   H������������#       H���   u+ƃ�    L��  H����  1�Hǃ       ��@  H�BH��   � ƃ   ����ƃ�    L��  ��   H����  � �   ��@  ����H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�BH��   � ƃ   �����ƃ�    L��  ��   H����  � �   ��@  ����L�ED��H���%  A�   H��H���	 ����������H�P�z�6���H�R�:>�)���H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �(ƃ  (H�E�����L�ED��H���P  �|$P H��(  �G����@���H�@H���D���D�����H�E�8�����H�U�:)HD������H��H��謔��H��u�D  H�x tH�@A��H��t�8/t�H�t$@H���	 H��H���x�  1�H����H��H��H��H�������H��   H��&H��H��H��H��   H9�@�,@��  �z���H=�   �.uϺ�   ƃ�    L��  H����  �   1҃�@  �H���	 A�   H������H� tfI��D��H���B  H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   � ƃ   I��D��H���  H�������I��D��H����  ����I�@�8)t
ǃ0     M�@D��H���  ����D��H����  ����L�ED��H���z  M��D��H���  �>���L9��������   ����<_�
���H�$       �   �   ��u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   @�4@��  L�������D��h  ǃ0     ����H��   �   u.ƃ�    L��  ��   H����  Hǃ       ��@  H��   H�PH��   �-ƃ  -L�E����H�	�	 A�   H�������.���E���n����a���M��D��H���  �^���fD  VSH��8M��H��L��toA�@��f��4  ��   X����L�D$ A�@H��H  ��4  H��H�D$(H�D$ H��H  �s���H�D$(H��H  �k��4  H��8[^�D  ǆ0     H��8[^�D  f.�     AUATUWVSH��(A� ��H�ˉՃ�LL���}  H�R�	 Hc�H�����  (tLH��   H�PH=�   u'��   Ɓ�    L��  ��  �   1���@  H��   � ƃ   L�F��H�ٿ:   H�5��	 H�n����H��   �*�H��H��H��H��   H9�@�<@��  ��  �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � M�@��H��H��([^_]A\A]�6���fD  H��   �   �?  H��   H�BH��   � ƃ   ��  H��   �   �l  H��   H�BH��   � ƃ   �  f.�     H��   �   ��  H��   H�PH��   � ƃ   L�F�=���f�     ����  H��   �   u+Ɓ�    L��  ��   ��  Hǃ       ��@  H��   H�PH��   �*ƃ  *�L%         H�=(�	 H��   A�    L�o	�- H��H��I9�H��   D�$D��  ��  D�'H��H=�   uκ�   ƃ�    L��  H����  �   1҃�@  �f�H�5��	 H��   �c   H�n�0�    H��H��H��H��   H9�@�<@��  ��   �>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �&ƃ  &H��([^_]A\A]�@ H�5��	 H��   �i   H�n	�,�    H��H��H9�H��   @�<@��  t��>H��H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  ��    H�5��	 H��   �    H�n�0�    H��H��H9�H��   @�<@��  �-����>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � H�5|�	 H��   �    H�n�0�    H��H��H9�H��   @�<@��  ������>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � H�5�	 H��   �    H�n�0�    H��H��H��H��   H9�@�<@��  �)����>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � H��   H�5��	 �&   H�n�0�    H��H��H��H��   H9�@�<@��  ������>H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � H�=�	 H��   A�    L�o&       �0fD  H��H��I9�H��   D�$D��  �N  D�'H��H=�   uκ�   ƃ�    L��  H����  �   1҃�@  �f�H�=��	 H��   A�    L�o�0fD  H��H��H��H��   L9�D�$D��  ��   D�'H=�   uκ�   ƃ�    L��  H����  �   1҃�@  �f�H�5�	 H��   �    H�n�0�    H��H��H9�H��   @�<@��  �-����>H��H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � I���l����     L�FM�������H�PH=�   u.L��  ��   ƃ�    H����  L�F�   1���@  H��   �(ƃ  (��H���M���H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �)ƃ  )H��([^_]A\A]ÐL�F�f.�     Ɓ�    L��  ��   ��  Hǃ       ��@  ����Ɓ�    L��  ��   ��  Hǃ       ��@  �����Ɓ�    L��  ��   ��  Hǃ       ��@  �d���ATUWVSH�� M��H�ˉ�L��L��tNA�I��uFL��A�   �
 �P��u1H�P�
����wL��H����1 ��  ���0  H� H��u�L��(  ��E1�I��Hǃ(      H���v  H��   H���   twH�BH��   �(ƃ  (L�E M��t��H������H��   H=�   ��   H�PH��   A�   I�����)H��ƃ  )�  L��(  H�� [^_]A\�L��  ƃ�    �'       �   H����  �(��@  ƃ  (Hǃ      L�E M���c����   �v�����   ƃ�    L��  H����  �   1���@  �K������  H��   �у����(��   H=�   ��   H�PH��   E1�I�����(H��L��(  ƃ  (Hǃ(      �  H��   H=�   ��   H�PH��   �)ƃ  )�s���f���  H��   �� �u���H=�   tTH�PH��   � H��H=�   ƃ   �T�����   ƃ�    L��  H����  �   1���@  �)���ƃ�    L��  ��   H����  � �   ��@  �������   ƃ�    L��  H����  �)�   ��@  ���� f.�     AVAUATUWVSH��@M��H��A��L��D����   ��0  ����   I�      A�   �_L��H��L��uBH�S��)�C   H��   H��   ��   ��*te����   D��H���g���H��   H�H��t[��0  ��uQ�C��u�L�C��A� u��H��3v�H�S��*�C   H��   H��   u�L�I��D��H���T  H��   H��@[^_]A\A]A^�L�I��D��H�������H��   H��@[^_]A\A]A^�M�@D��H��H��(  Hǆ(      ����A��H��   H��(  ��   H�PH=�   u*��   Ɔ�    L��  H����  �   1���@  H��   �.Ɔ  .H�CH�h�E ��F��   ����3w/H�      H��s�   H�m�M ����3wH��H��H��u�I��D��H���L���H��   H��@[^_]A\A]A(       ^�H�--�	 A�:   L�u�. H��H��H��H��   I9�D�,D��  �U���D�m H=�   uͺ�   Ɔ�    L��  H����  �   1҃�@  �H���	 H��   A�{   L�s�&H��H��I9�H��   D�,D��  t<D�+H��H=�   uҺ�   Ɔ�    L��  H����  �   1҃�@  뭋EH�\$ H�M�	 H��D�@���  H�ڋ
H����������!�%����t�������  D�H�JHDщ� �H��   H��H)�t`L�,�"H��H��H��H��   I9�D�4D��  t8H=�   D�3uҺ�   Ɔ�    L��  H����  �   1҃�@  �H���	 A�}   L�s�&H��H��H��H��   I9�D�,D��  t8D�+H=�   uҺ�   Ɔ�    L��  H����  �   1҃�@  �H�m�E ����fD  AVAUATUWVSH�� M��H�ˉ�M��M��L��t#�P���$  H� H��u�E1�M���H���|���H��   H=�   �  H�PH��   � ƃ   H���   t]H�BH��   �[ƃ  [M�$M��t��H���q���H��   H=�   trH�PH��   �]ƃ  ]H�� [^_]A\A]A^�L��  ƃ�    ��   H����  �[��@  ƃ  [Hǃ      M�$M���}����   돐��   ƃ�    L��  H����  �   1���@  �c����H�@�8*uL��E1�M��H���W���H��   �������   ƃ�    L��  H����  � �   ��@  �����H�5��	 H��   �    L�v�'f�H��H��H��H�� )         I9�@�<@��  t>�>H=�   uӺ�   ƃ�    L��  H����  �   1҃�@  ��    E1ɉ�M��H������H��   H���   t H�BH��   �)ƃ  )�����D  ƃ�    L��  ��   H����  �)�   ��@  �����UWVSH��(A�81H��tH��([^_]�b���f�I�@HchH�pH��toH��   H��% H��H��H��H��   H9�@�<@��  t>H=�   �>uӺ�   ƃ�    L��  H����  �   1҃�@  ��    H��([^_]��    WVSH�� A� ��0H�ˉ�L����   H��   H�PH=�   ��   H��   I����H���(ƃ  (����H��   H�PH=�   u*��   ƃ�    L��  H����  �   1���@  H��   �)ƃ  )H�� [^_��     H�C      H���W�����H�� [^_�������   ƃ�    L��  H����  �   1���@  �1���D  f.�     AWAVAUATUWVSH��(I�@��H�1�H�ˀ:f�}  I�E1�L�xL�`A�?;�A  ��<  ǃ<  �����B<R�^  �T  <l�'  <r�(  H��   H�PH=�   ��  H��   M����H���(H�5v�	 ƃ  (�B���M����H������L�fH��   �.   �, H��H��H��H��   L9�@�,@��  ��   �.H=�   uϺ�   ƃ�    L��  H����  �   1҃�@  � M����H������M����H������H��   H�PH=�   u*��   ƃ�    L��  H���� *        �   1���@  H��   �)ƃ  )��<  �   H��([^_]A\A]A^A_�<Lu�H��   �   ��  H��   M��H��A�.   H�5��	 L�~H�PH��   ���(ƃ  (�����M����H���.���H��   �/D  H��H��H��H��   I9�D�,D��  �����D�.H=�   uκ�   ƃ�    L��  H����  �   1҃�@  �f�M�wM����� H�5|�	 H��   A�(   L�v�,fD  H��H��H��H��   I9�D�,D��  t>D�.H=�   uҺ�   ƃ�    L��  H����  �   1҃�@  �fD  M����H���#���M��������   ƃ�    L��  H����  �   1���@  �4���ƃ�    L��  ��   H����  Hǃ       ��@  �C���f�     UAWAVAUATWVSH��  H��$�   D�1A��_H��I��M���~  H�=T�	 H�޹   ��� 1���u2�C��$<;w'H�     H��s�C	<D�{  <I�s   H���8�  H�]�H���E�   H�H�]�D�H�E�Ic�D�E�H�@�E�    H���U��E�    H�E�    H�E�    �E     �^  H)�Hc�H�|$'H��   H��L�<�    H����6  H)ă�L�}�H�D$ H�E��=  ����   ����   �{_L�sL�u��~  L��D�E��n�  D�E�E����  ���E�   ��       ��  ��        H�]�L�4�   ��   1҃�H����M��E1Ƀ�C� n��H�]�H��H����  H�H��H�]��u*f�1��p  f�     +       H�M������H��H�E�� H��t؄�u�H�}I��Hǅ      H��H��\  ƅ   H��l  L��   L��(  Hǅ0      Hǅ8      Hǅ@      HǅH      ǅP      HǅX      Hǅ`      Hǅh      Hǅp      Hǅx      ��m����|  �   Hǅ�      Hc�l  �Ѕ�HN�H����|  �e  H)ą҉�O�L�D$ H�H���K  �   H)�L��`  H��I��H�D$ H��p  ����H��  H��H��L��(  �D ��   ��@  1�����H���  [^_A\A]A^A_]�D  A��_�f����{Z�\���H���   H�]�H�]�H��蓚���E�H����   H�E�� �M���f.�     �yZ�   �s��������{Z�x���H��1�H�]�H�]�H���<���I������@ 1��{
_�����1�<I@�ƃ��t���@ H�]�E1��{���@ H�EȋU�L)�;U���   Hcʃ���L�IH�M�N��A�A    �U���   I�    M�AA�AI��M   H���Yk��H��L�E�A� <.�i���A�@�P���vi<_te��0<	��   A�L�� ��.�g����x�WЀ�	�W����PH�H�B�<	w�     H����B�<	v�H���E1��l���D  A�PI�@�J���wH����J���v��_t��A� �����ATUWVSH��@H��H��L��L����   H��t	M����   L�D$ H�D$     H��s���D$8    H�D$(    H�D$0    �r�������   �D$8H�\$ ��t]H��A�   ��   H����   H�����  H;E swL�@H��H���X�  ,       H��H����  H��t�    H��H��@[^_]A\�@ H��L�d$0u�H��tI��uZ�����1��ϐH��t�����1�H��H��@[^_]A\�D  H���H�  L�e �f�H��u��f�     H�L$ �&�  H��t������1��r���H��u�1�먐f.�     H��(H��tH��t�]���������H��(ø���������������H��(H�eb	 H� H��t��H�Tb	 H�PH�@H�Eb	 H��u�H��(Ðf.�     VSH��(H���	 H������t9��t ��H��H)�H�t��@ �H��H9�u�H�~���H��([^��f�� 1����D�@J�<� L��u��f.�     ��! ��t�D  ��!    �q����H�%-H ���������1�Ð������������ATUWVSH��0H��	 H�2��-�+  H9�H�D$     tH��H��	 H��0[^_]A\�f�H�L$ �IF H�t$ �F A���F ���EF H�L$(���pF H3t$(D��H�������  H1���H1Ɖ�H1�H!�H9�t%H��H��H���	 H���	 H��0[^_]A\�fD  H��] �f���H�3��-�+  ��f.�     UVSH��H��pH��H��  �"F H��! H�U�E1�H���F H����   H�U�I��I��H�D$8    H��  H�T$0H�U�H�L$ 1�H�T$(H�U���E H��! 1�H�5! H�v% H�	 �   H�U% H���	 H�E�H���	 H�E���E H���	 � F ��D �	 �H����E �{�  H�EH� ! H�EH��  �{�����������H��(��t��t�   H��(�f�     ��  �   H��(ÐVSH��(H�#�	 �8-       t�    ��t��t@�   H��([^�f�H��_ H�5�_ H9�t�H�H��t��H��H9�u�   H��([^��Y  �   H��([^� f.�     1�Ð������������H��XH��$ H��t,��$�   �L$ H�L$ H�T$(�T$0�\$8�D$@�АH��X�D  f.�     H��$ 鼽  @ VSH��x)t$@)|$PD)D$`�9��   �H���	 Hc�H���H���	 H�q�DA �y�q�   蚽  �DD$0I��I���|$(H�x�	 H���t$ 肼  �(t$@1�(|$PD(D$`H��x[^��     H�h�	 ��    H�y�	 �|���@ H���	 �l���@ H���	 �\���@ H�i�	 �L���@ H���	 �<���������Ð������������H���f�f.�     H��Ð�����������ATUWVSH��PHc5s# ��H��H��L���f  H�_# 1�H���H�H9�rL�@E�@L�H9���   ��H��(9�u�H���A  H��I���R  H�# H�4�H��H�L�` �     �D  A�L$H�T$ A�0   H�H��" H�L0��B H����   �D$D�P����t��@��ub��" ��s)@����   ��t�E @�����   H��P[^_]A\É���H�T���H�T�r���1���H�L 9�H�r���H5Q" A�@   H�L$ H�T$8I��H�NH�V�$B ���n�����@ H��	 ���lZ	 �E ����D=��D;��p���1���������D=�f�D;��X���H��! H���	 A�T$L�D0�#Z	 H�\�	 H���Z	 � UAWAVAUATWVSH��8H��$�   .       ��! ��tH�e�[^_A\A]A^A_]��s!    �  H�H��H��   H����7  L�% �	 �J!     H�5��	 H)�H�D$ H�8! L��H)�H��~�H�����   ����   L9��y���L�vI��L�-��	 H�}�M)�I��N�d��
fD  I���NA�   H���L��L��E��>���M9�uً�  1�L�%�@ ������f�H��  H�D� E��tH�PI��H�HA�ԃ�H��(;w  |�������N���Q����V��u�VH�� ���8����F���-����V���/  L�-*�	 H��I�    ����L�u�L9�rH������   �� �   ��@��   H�A�   L��H)�L�H�U�L���X���H��L9������N��VL�L��L�u�D�L��L��M��I��  ��fE��MH�I)�M�L�E�A�   ����멐�L��I��L	�E��II�A�   H)�L�H�U�L��������y������u5D�L��L��M��I�� ���E��MH�I)�M�L�E�A�   �����>���H�g�	 H�E�    �bW	 H��	 �VW	 ������H��(�=�  �wc=�  �s{=  ��  ��   =  ���   =  ���   1ҹ   �9�  H���/  H���<  �   ��1�H��(��     =�  ���   w7=�  ���   =�  �uo1ҹ   ��  H��toH��tX�   ��1�H��(�=�  �ti=�  �u<1ҹ   貵  H����   H����   �   ��1�H��(Ð=  �t�=�  �t&�   H��(��     �   �   �a�  ����1�H��(�D  1ҹ   �D�  H���[����   �   /       �+�  1�����@ �   �   ��  1������f.�     �   �   ��  1�������   �����ATUWVSH�� �  H�ŋ` ��u%H��t H���	 �F    �  H��t�   H�� [^_]A\�@ H�9 �0   1�H�+ H���H�L�%�����    H���H�I)�H���.�	H��H��D�g�H�K�HH��H��H)�C��K�H�� t2H���u  H��u�H�����q���D  H�� I����; �W����    ��@ SH�� H��H�ˉ������ ��CCG ��   =�  �wh=�  �s|=  ���   ��   =  ���   =  �u1ҹ   蒳  H���Q  H���  H� H���  H��H�� [H��@ =�  ���   wX=�  �tF=�  �u�1ҹ   �9�  H����   H��t��   �и����H�� [��     �B�7��������H�� [�=�  �t�=�  ��j���1ҹ   �ݲ  H����   H���K����   �и�����=  �t�=�  ��+�����     1ҹ   蔲  H���[����   �   �{�  ������S�����   �и�����A���1��:����     �   �   �A�  ������1����   �   �(�  ��������   �   ��  �����������������UWVSH��(H�A ��8 H� H��t3H�-$: H�=9 ����H���ׅ�uH��t	H�CH����H�[H��u�H�� H��([^_]H�%"9 fD  UWVSH��(�� 1�����H��u��H��([^_]ú   �   �M�  H��H��t=�(H�� H�x�N8 H�k H�0       � H�] H�C��8 ��H��([^_]þ����뚐SH�� �= ����u1�H�� [��    H�9 ��7 H� H��t�9�u�O�9�t)H��H�HH��u�H� �<8 1�H�� [��     H�QH�P�3�  H�� �8 ��@ H�PH��H�� ��SH�� ����   r0��t��u�� ��t�G����
D  ������   H�� [Ëb ����   �T ��u�H�@ H��tH�Y袰  H��H��u�H�C H�     �     ��6 �fD  � ��t��    �   H�� [ÐH�� �7 �ې�����t���������HcA<H�1��9PE  t�1�f�y���f�f�9MZt	1��fD  ��@ f.�     HcA<H��AH�D�I��t)��H��L�L�(D�@I9�L��wHH9�wH��(L9�u�1��f�f.�     WVSH�� H�����  H��wkH�T�	 f�:MZu]H���E�����tQHcJ<H��AH�\�A��t9��H��H�|�(�	H��(H9�t"A�   H��H���Y�  ��u�H��H�� [^_�f�1�H��H�� [^_� H��(L���	 fA�8MZH��uWL���������tKIc@<H��L)�I�A�PA�@��I�D t+��H��L�L�(f�D�@L9�L��rPH9�rH��(L9�u�1�H��(�f�f.�     H��(H�U�	 E1�f�:MZtD��H��(� H���8�����t�HcB<D�DD��H��(�f�H��(L��	 fA�8MZH��uRL��������tFIcH<L��AH�D�I��t.��H��H�L�(f.�     �@' t	H��tH��H��(H9�u�1�H��(Ð1       H��(H���	 f�:MZuH���������    HE�H��(�fD  1�H��(�f�     H��(L�e�	 1�fA�8MZH��tH��(� L���H�����t�Ic@<H��L)�I�A�PA�@��I�D t1��H��L�L�(�     D�@L9�L��rPH9�rH��(L9�u�1�H��(Ë@$����H��(�D  f.�     H��(L���	 fA�;MZA��uXL��������tLIcC<L؋��   ��t;�HH�L�@��t*��H��H�D�(D�QL9�M��r	DAL9�rH��(H9�u�1�H��(�L�u��@ A��H���J��u�B��t�E���BL�H��(Ð���������QPH=   H�L$rH��   H�	 H-   H=   w�H)�H�	 XYÐ�������������H��81�A�   H�L$@L�L$@�CCG"��2 H�D$@�   H�P0I��H�D$     H�T$(L� �   �P�   H��8Ðf.�     H��(��wHc�H�D�H��(���  �@ H��(��wHc�L�D�H��(��ͫ  �@ H��f�f.�     H�AÐf.�     H�A�    �D  H�QÐf.�     H�A H�@8��    H�Q H�B� HBÐH��8E1�H�T$(�B2 H��t� HD$(H��8�1�H��8�fD  1�� f.�     H�A H�@��    AUATUWVSH��h�A� H��H��M��L����   �H�y ��CCG!��   I�I(��CCG"L�L$PH���   H�L$0I�	H�L$8�ﾭ�H�L$@H�L$H��   ��CCG uv�L���   H�t$0�   H�t$ I���   ��$�   ��tH���)  H�D$8H�k(L�K A�   �   �CCG!H�C0H�D$HH�C8�2       �0 ��   H;i(��   �   H��h[^_]A\A]� I�A(H�Q8H���   ��H�G0H�t$0�
   I��H�t$ �   H�D$(L��WL��
   �F���L�l$0I���   L�l$ �   ��$�   ��t���uiL�l$ I��L��   �   ��$�   ��uHH�D$HH�oI��H��H�T$8L�L$@H�G(H�W H�C8H�F@�C   H�k(H�S0H�D$(L�d$ �70 �>�  I�A@I��H�Q0L�D$ I��H��H�D$(�0 ��  �D  f.�     WH�� 1�A�   H�L$0L�L$0H�ʹ   H��H��1��H��CCG ��/ �   H�� _�D  f.�     UWVSH��  1�H�T$8H�˹   Ǆ$�    H��$�   H���H��   H��H�\$P�H�H�l$0H�CCG    �D$H   H�D$0H�CH��$�  H��H�D$XH�C H�D$`H�C(H�D$h�/ H�S I��I��H�KH�t$(H�|$ �/ �
�  ��H��(H�y u
�������  ������@ H�A    H�A     H�A(    H�A8    H�QL�A0�S��� H�AH��tH�ʹ   H��Ðf.�     AWAVAUATUWVSH��x  1�H��$�   I�Ϲ   H�D$@    H�\$pH��I��H�D$H    �H��
   H��H�D$P    �H�L�l$@H�D$X    H��$�  H�D$`    Ǆ$�    H����- H�\$`H��$�  H��$�   L�%�- H��$�   H�=�- �Z�    H�CH�S1�H�D$8    H�D$0H�C8L��$�  H�D$(H�l$ ��L��L��H�C0A�ׅ�uOH��$�  H��t$H�\$`H�H�SI��A��H�CH�\$`L�KM��u��   H��x  [^_]A\A]A^A_�D  3       �   �����������WVSH�� H�9H��H��t1�H�D�H��t	H�H�蹥  H��H9�u�H��H�� [^_顥  �H��(H�� 1���  H�����H�� ��  ��uH��(��ť  �f�f.�     ATUWVSH�� H�qH��H��t=�T ���  H��H��tgH�(H9���   H��L�M���   L��H�� [^_]A\�H�f���H�� ���  H� �~�  H�wH���  H�� ��  � H�N!�   ��  H�n H��H���  �� H�(H����  �q���H�wH�/H����   H�L5�9�  H����   L�L0H��I!�I�A�H�WI��H����   L����  I��L��+���fD  L�d- H��H�F L9�LG�J��   蘣  H��H��tzL� H�L�I)�1�N��    莣  � H�����  �����H�M蚣  H��t?H� L�H�h����H�� H�pH�5� H�w�����D  L��1��6�  I���P�����  ��     H9sH�H�A    L9AsL�AM��tH9t�L�IÐ�����SH��@L�DE	 H�D$8H�D$ L�L$4��  ����w+H���	 Hc�H���fD  �\$<�T$8��  �H�� H	ӨtH�؉�H��    �H�� H	�fHn�H��@[��    H�      ���@ 1����L$4�T$<��3  ��������	�H�� H�ڋ\$8H	�� �\$<H�� H�ڋ\$8H	��H�      ��r����������������H��HL�uD	 H�D$8H�D$ L�L$<��  ����wwH�б	 Hc�H����    �  ��с�   ��E�fn�H��H�D  �T$8��f.�     �L$<��� 4         �L$8������ 	��D  �  ��f�     1�롐�����������H��H��������t=�L$=f�D$>謢  H�T$>A�   �D$(   H�T$ L�D$=�   ���n( �D$>H��H�VSH��X1�H��H��H����   M���0  �A�	A�    �҉L$L��   ��$�   ��   ����   L�L$8��$�   L�D$0��' ��tfL�D$0L�L$8I����   H�t$ A�   I���D$(   �   ��$�   ��' ����   �   H��X[^�fD  1�f�H��X[^�@ ��$�   ��u5�f��   H��X[^� �T$MA�   �D$(   L�D$LH�t$ �f��D$(   A�   I�غ   H�t$ ��$�   �,' ��t�   �m���f.�     ������Y����Ѡ  � *   ������D����A�������4����UWVSH��X1�H��H��f�D$NL��H�D$NH��L�D$8HD��   ���à  L�D$8H��H��L��
 �l$(H��LEΉD$ �%���H�H��X[^_]�f.�     AVAUATUWVSH��@H��
 M��L��I��HD�H��L���[�  1�A���I�  M��A��tZI�H��tRH��tdH��u�FI�H�H��H�H�H9�I�v/I��D�d$(I��H��I)�D�l$ �������H9�v��uI�    H��H��@[^_]A\A]A^�D  H�t$>1�D��f�D$>�I�H�H�H�I�D�d$(I��I��H��D�l$ �)������� UWVSH��H1�H��H��L��f�D$>�s�  ���t�  H�ۉl$(I��H�{	 �D$ HD�H��H�L$>I�������H�H��H[^_]Ð�������UAWAVAUATWVSH���   H��$�   H��H���   �Ɲ  H��H� 5       � �E��%�  I�ƍ@�E�H�H��H�������H)�I��L�d$0�I��A�D��)�A��苝  ��u�D�E؉�E���(  I�GE��E�,$I�T$t#A�NM�D�H���H�H���ɈJ�tI9�u�� A�$<-��   1�L��<+f�U�I�T$HD�A�   H��H��	 誝  ��uvL�vA�   H��H�լ	 L��艝  H�M�H�E�    H���   ���A    LD�1�f�A��  f�E��E�f�E��9  M)�F�,7D��H�eX[^_A\A]A^A_]�f�H�s�	 A�   H����  ��uJH���   H�M�H��   �  H�E�    H�E��E�L�vf�E��E9  � I�t$�����f�M�����1�H�E�    f�E �H�E�    <0�$  H���<0t��E�   L�EE1�1҉}�H�M�L�e�L��E1��E�    E1�A��E��H�M�L�u�]��% �U�f��tG	]�A��A�� A	�A��H����؃�0��	v�8E��:  E���  A�   ��f�     H�E�A��A���1�L�HL�Pf.�     A�A��A��f��AH��A��A����AE�I���fA�AM9�u�L�M�1�1�L�U�f�E 1�L�ML�OL�U�A�A��A��f��AH��A��A����AE�I���fA�AM9�u�H�O�     �A��A��f��AH��A��A����AE�H���f�AL9�u�H�U�H��D�E��`3  H�U�1�H��H�    H�G    f�Gf�]�;3  D�E�����f�DE����E��D�m�<E�]ȋ}�L�e�E����  D)ۅ��$  f�}� �  L�uH�u�foE�L�}L��L�u�)EL�N1�1�f�M 1��A��ʃ�f��H����6       ����E�I���fA�AM9�u�L�N1�f�     A��ʃ�f��H������E�I���fA�AM9�u�L��H���Y2  L�N1� A��ʃ�f��H������E�I���fA�AM9�u�f�} u&foE1҃�f�U )E���   f��f������H�u�H�M��8  ��P�5  H�E�H�E�    H�@
    �E�H���   H�M�f�E���5  �E̅�t(H���   �(���}���������zt9H�E�f%�f=�tE�������I�������D  H�E�H��H�� �����	�u��f�  � "   ��DE�E��D�m̋]ȋ}�L�e�E���$����L������E���c  1�����H�M�H�u��7  ��P�!����U�A�N@  E1��D$(P   H�M�A)��D$ @   �J9  �E�E�D�M�E1����D$(@   H�M��D$ @   �!9  ������U�A�N@  E1��D$(P   H�M�A)��D$ @   ��8  �E��E�   �E�H�E0H�E�H�'�	 L�=�	 H�u���L�uM��d���H�E��	 �E�   ���f�     I���M9�t��t�M��L��L��L�M��?<  L�M���H�U�L��H�u��/  �}����   H�U�H�M�D�u2Du���2  ��A������E�������E�    ������F<-�9  L�v�   <+u	A�FI���PЀ�	�������q  ���\P�I��A��PЀ�	v����N  ��q  L���J���D�]�E1�H�E�    H�E�    fD�U E���_  �E�A��  L��H���   fD�M�H�M�f�E��,3  �Y����E2D�u�H�U�H�M�A)��o/  ��A���?  �E�����H�M��5  ��P������U�A�N@  E1�7       �D$(P   H�M�A)��D$ @   �7  �E�ۉE�������� ���|(H�E0���E�����H�E��	���L�v�F���������L�}0H�z�	 L��L�}��n-  �E2L��D�u�H�U�A)��.  A���?  �E������Eи ���)؉�������q  ~ZH�M�H�E�    �E�H���   H�A
    f�E��2  D�E�E���N���L���%����E�H���   H�M�f�E���1  �)�����L������f�f.�     WVSH��0H��L��H��H�D$     H�T$ H��H�D$(    ����H��tH�H�H��l$ H���>H��0[^_Ð��H��XE��D��f�T$huf��� wR��   H��X�H�T$LD�L$(A�   H�T$8L�D$h1�H�L$ ���D$L    H�D$0    �. ��t�T$L��t���  � *   �����H��XÐWVSH��0H��H�ˉ�H�D$+HD���  ����  ��A��H��A���K���H�H��0[^_ÐAVAUATUWVSH��01�I��I��M���ʔ  ��軔  I�] ��H��tM��tkM��u>fD  I�] H��H��0[^_]A\A]A^�f.�     H�I�H�A�~� tqH��I9�v��A��A��L���������H�������f.�     L�d$+1���    HcЃ�H�Hր|+ t/H���A��A��L���i������� I�E     H���S���H���J���������H��Xf�L$J�D$L    �ғ  H�T$LA�   H�D$0    H�T$8H�T$I��H�T$ L�D$J1��D$(   �| ��t�D$L��u�D$IH��X�f.�     ������ꐐ�������WVSH�� H�5R�	 1�H�٢	 H���@ H�H��H��聑  ��t����u�1�H�� [^_�H�8       �	 Hc�H���DH�� [^_��#�  �����������WVSH�� 1�H�ˋIH�s�ʃ���tH�3�C    H�� [^_Ð��%  t�H�;1�H)�H��~�H���J�  A��H������  H�H9�u�SH�s��%�   t����1��S롃K �����H�s�D  WVSH��0A��H��H��t-A��tGE��ulH�T$(H�t$(H��H���%�  H��0[^_�D  H�t$(H���C�  ��u2H|$(���     �3�  H�t$(H��薑  ��藑  H�H�|$(른�����葑  �    ������@ AWAVAUATUWVSH��(H���h�  H���     �B�  �ǋC��y�C    1�A�   ����  H��H����  �S��  ��   H�H�CI��I)���un���  L��H����   ���   HcC����   L�=�	 N�$A��A��A��A��Mc�I��I�J��B�|( ��   L)�H��pf�     L�ɵ	 A��L��A��Mc�M�A��A��I��O�A�x �m���H9��a���fD  E1��8
A��H��L�H9�u��C���D  HcCH)�H��H��([^_]A\A]A^A_�D  H����E1�H����֏  I��   w�S�   ��  ��tHcC$I�J��B�D*tH��H)��     H��1�A�   ��脏  H9�u�H�SN�"L9�sf.�     1ɀ:
��H��I�I9�u��C u"L)�H�4(�A���f.�     H�������+���M�L$L)�H�4(�����N�  H�������    ����f�f.�     WVSH�� H��H��D����  H���     tr��wm�c��tUH���J����C��t3����CH���͎  A��H�9       ���蠎  H���������H�� [^_�@ %	  ��	u��C$   ��H��1��#���H��虎  �    �������f�f.�     VSH��(1ۉ�詎  H�^�	 �0H�J��   �H���<��t#��9�u��G�  H�0�	 �T��H��([^� �F��v8��   ��v��  �    H��([^���  �    H��([^�f�     ��  �    H��([^Ð�������������H��8H�T$(�2�  ��uH�D$(H��8�@ H�������������c�  �����������VSH��8H��H��t2H�Z�L�L$ H��M��1�A���9M  ��9�O�Hc�� H��8[^�@ L�L$ H��M��1�E1��M  H��8[^Ð���VSH��(LcIH�AH��M��J���fD  H���@�    H9�v ����t���H��H��([^�f.�     D;C}A��H��D�CB�D�   H��([^ËC�H�d}  H�SH�HH��HcCL��   �x�  H��H���=~  LcNM���@ AWAVAUATUWVSH��H�H��L��M��H�T$<L�D$8�ą  �T$8D�.H�ËD$<D)�Ѕ҉T$8�D$<��   A��5��   ��$�   ��  ��$�   ��  H����  �T$8H�ى���u  H�������    H��D��K��)�EQ�Hc��T���9��o  ��u�{���   H��A�    �u  �D$<���D$<�VD  ��$�   E1���t
�~�k  H��� }  D��H��H[^_]A\A]A^A_�D��$�   E1�E��t�1�E1����_  �V9���   A�щT$<A)�E9�|uD�vE��ulA�q���~����  ���$�   t����   ����H��Hcҋt�D:       ��!���t  H��$�   ���    ��  ���P   �D$<DE��"�     H��$�   �C    E1�� P   �ЉE I��D��L���5�  H��$�   A�   D	8������V9�}�H��$�   ��E1��T$<� �   �K�  � "   �D$<�C    ��     �Ѓ�ui��$�   E1���������C����H����  �T$8H�م�����   ��s  E1��D$<���� H�����  H�ËD$<����f.�     ����HcɋL��������H��賆  ������   �T$8H��A�   �s  �D$<�?�����H��D�L$,��  D�L$,���W��� �[s  A�   � �D$<A�    ����H��A�`   ����H�ËD$<����H���/�  �T$8H�م���u��s  E1��2����T$8H����f�f.�     HcQH�AH���f�H���@�����H9�v���t����@ SH��0�ZH����9Y|bL�@������t?���HHc�I��L9�vI��A�@�����L9�w��t�    )�A�h�H��0[��    �HHc�I��L9�w�H��0[ÉT$,��y  ����x  �T$,�D  AWAVAUATUWVSH���   )�$�   )�$�   D)�$�   H��H��$H  L��$P  L��$X  ��  L� L���I�  H��Ǆ$�       I��H��$P  HǄ$�       H��$�   H�!�	 HǄ$�       D�� A��-�D$@�E  A��Hc�H����     H��$H   �   Ǆ$�      tH��$H  H�(��$�   (�$�   (�$�   D(�$�   H���   [^_]A\A]A^A_�fD  �D$X    H�rH��$�   D�BE��t�A�;       �0�D$D    ��   H��$P  H��    �    �@�D$tA���PЃ�	�    v1��   D��B�|@�H����H��$�   �D�H�A��A��	��   ��~σ�Ӎ��TP����D$X   �Z���f�H��H��$�   D�A��-�����fD  A��0H���D$X    �D$D    �C����F<X��  <x��  H�FH��H��$�   D� H�@A��0t�E����  �D$D   �����E8$�r  A��1��D$P    E1�A��A���A��E��   E1�E����  �|$D	���  E����  ��Nt��  ��i�  ��n��  H��$�   H�ݗ	 H��輁  ����  H��$P  Ǆ$�      H��$X  L��$�   �@�D$D���H��$�   �8(��  L��$`  H��H��$P  ��p  ��$�   H��$P  H��$X  L��$�   �@����P  D��	�D$D�!  H��$�   H�EH��$�   �E<+�  E1�<-uA�   H�EH��$�   �ED�@�A��	��  ��0u&H��$�   L�@D  L��$�   A� I����0t�D�H�E1�A�������L��$�   D�@�M�kL�\$HL��$�   A�CD�H�A��	w5M�Kf.�     G��L��$�   M��I��F�D@�A�A�D�X�A��	v�L+l$HI���q  A��N  �d  E��A��E��EE��������I�C  f�L��$�   H��$�   Ǆ$�      D  H��$H   tH��$�   H��$H  H��D$X��t��$�   M�������H��$`  �T$@��  H��$�   ��t  �����H��$X  H�A    �|$\�8�D$t����  �P   ��@��$�<          ���  � "   L��$�   �]���Ǆ$�      D�\$XH��$P  D+D$P�@D�D$p�D$D����D)ك��L$dtA�K���L$dt�������D$d��f���۽   �H*�AD�A��AN�A��	��$�   ~'H��	 �E�f���H*�H��Y��X���$�   �|$@5�{  A���q  �|$p ��  �  �D$p���^  ��$�   Lc�H�B�	 B������  �ʺ5   )�H�e�	 ���$�   ��5D�T$d�����BY��D$ L��$�   H��$�   L�D$0D�T$(��$�   L��$`  L��$X  H��$P  ������������1��    E�D$E���F  D:A�u���H��I���H��I��E8�Z���E�$I��E��u��L��$�   A� �\  D�@�1�A���D$P    A��	��  E��E��L��$�   �A��  ��I�AH��$�   A�AD�@�A��	v��H  �    �D$pD��)��Ń� ��  ���t H��	 H���$�   �Y���$�   �����  ��$�   H��$�   L��$�   �y  ��$�   D�|$@H��$�   �$�   A��E)�E�퉬$�   ~'D��H���j  ��$�   D��D��$�   D퉬$�   �*+D$@����$�   H��$P  �@�D$D��9���  H��$P  �@9��D$\��  )Ń� �L  ��  �D$t�T$\����$�   �?  ��$�   ��9��-  H��$�   H��$X  H�A    � �A    Ǆ$�   P   �I  L��$�   � "   ����fD  �D$XH��$�   L��$X  L��$�   H��$P  �D$ ��_  ��=       ��$�   �	���H��$�   L��$�   H��$H   �����H��$H  H�(�r���@ H��$�   E1������������`  H�{�	 D�P�E1�E��A���J �     ��$�   ���с������  �?����$�   ���  A9���$�   A������Y�A����$�   u�D�Ѓ���$�   A�Ё����A����  �?A���  ����$�   ��$�   B����������H�Ģ	 f(�1ɨt	�Y
�   H����u���`�����$�   f(��N�����0�k  I��1�L��$�   A� ��I����0t�D�@�A����  �D$P    E1�A�   ����@ H��$�   ���s  �$�   H��$�   ����H��$�   �D$    H�D$0�D$dH��$�   �D$(���� ������݉��t H���	 H���$�   �^���$�   ����n�����������  H�c�	 D�P�E1�E��A���J ��$�   ���с������  �?����$�   ���  A9���$�   A������Y�A����$�   u�D�Ѓ���$�   A�Ё����A����  �?A���  ����$�   ��$�   B����������H���	 f(�1ɨt	�Y
�   H����u��+���@ �D$D    H��$�   Ǆ$�   �   �@    ��{  H��$X  � "   H��$P  �@���D�T$DL��$�   E������D�L$tL��E���$�����$�   A�H��0�����~�����c�����$�   �����fD  �D$\�D$D   ��$�   A����H��D�t$ E����u  �|$pH��H�D$h1��D~�	 ���څ�I�>       I�1�T$P�D$`H�FH�D$x�D$@�x����$�   ��$�   ��   D  �q  �L$DH��$�   ��uKA�T$��9P~Hc�H���L�A�T�����9�}"�T$\9�$�   �  ��$�   D�l$D@ L���l  L���l  ����  ��$�   �$�   ;D$Tu;D�l$HE��t1�Y5
�	 f(��\�	 f(�fAW�f.��h  f.��~  D�d$DE����  H���k  H���k  L���k  H���k  H�t$h�N�~j  H�T$xH�HH��HcFL��   �x  H��$�   �H�Qj  H��$�   H�HH��HcBH��L��   �]x  ��$�   �   D��$�   �4l  I���A)����  �D$PD�t$`D�,D�+\$@�L$\��$�   ��)�D)��9�O�A�\ A�D9�D��N�A9�ANŅ�~)�A)�A)ŋD$P��t-L�����!m  H��H��I����k  H��H�D$H�j  H�D$HH��)�� �$  �  �D$p��~�T$`H����l  H��E��~H��D���Fn  H��E��~L��D���3n  I��H��H���eo  �xH���h���  LckL��H���C    ��n  �T$d���/  ���'  �Ѓ���D1�D9��b  E����  �5Ë	 E1�Ǆ$�   !   �D$H    Ǆ$�       f(���$�   ��$�   �;D$@�T$T}�D$D�i  H��$�   f(�L��$�   � q  ��$�   I�ƅ��.  tH���Dm  I��L��$�   E��L��L��������
  �PH��$�   ��A9T$~ Hc�H���L�A�T�����9�������T$D���T  ��$�   ��;D$@��$�   �����D$D����?       ���]  ��  L��H���r  ���	 f.���  E����  1�A���D$D�=  �5q�	 �D$H    A�   Ǆ$�      f(�����H����El  H�������D�t$`D�l$PA)��4����   H���l  L��$�   H��$�   ��$�   ��g  L����g  H��$�   �9a  �D$D    ���/���f.�     Ǆ$�      �T$\9�$�   �*����T$@L��$�   ����  E�XE��������$�   �   A����H��E�T�E��������� Lc�9�u�A��~K�T�A�������A9ɉ�������$�   L������$�   �D$@��$�   ����H��$�   D  �l$D����  ��$�   H��$X  H����f  H����f  L����f  H�L$h��f  H����f  H��$P  ��$�   9x�V����@�D$P������  ����  �������H��$�   �f  H��$P  HǄ$�       H��$X  Ǆ$�      �@�H��$P  H��$`  ��A��H�H��H��H9�sH���@�����H9�w���������    )ȉ��j����� ��	 f(�A�����	 �Y�����A��A�ŉ�$�   E��f.���   �,�f���*��D$H�D$d���\���  ���F  E��u.f.=��	 v$�D$H�0   f���T$H+�$�   �*�$�   1�����f.�������I�	 �\�f.��������$�   	�$�   �����     ��H���f]  ������D�t$@H��$�   E��A)�D����h  D��$�   D)�$�   H��$�   �_����     f(��D$H@           1������5��	 �D$H    1�E1�Ǆ$�       f(������@ �   H����\  �D$H    ��$�   ��$�   �F���fD  ��H����\  �����f.������1�����E1������fD  ��$�   �D$D�D$@+D$D�� �D$D����H��$�   �T$D�   ��g  H��$�   ��$�   +D$D�D$D    ��$�   �����f��D$D    ����� E���'���1������T$p�����E���H�z�	 ����$�   H��^�H��$�   �D$     H�D$0�D$dH��$�   ��$�   �D$(�����L$p�%   D)�9ʉ������H��	 �   ��$�   D)�Hc��YʋL$p)�Hc��Y��H��$�   H���	 H���m  �������H���	 H��H��$�   �m  ��u	H��$�   Ǆ$�      ����L�A������H��$�   �҉�$�   ��  ��������H�      Ǆ$�      H�A�������������$�   �K���E����  Ǆ$�   !   A���-����L$\9�$�   �����D$D����H�ٺ   �f  L��H��H���g  �������Ǆ$�      �D$D    �D$@H��$�   )�$�   ��$�   �Z���H��$�   ����E����  D�D$DE���V  ��$�   L��$�   ��I�@��Hc�H��H9�s%A�x�I�@t�"  f�H���x���  H9�r�у�t������Ѓ���  H�      �L$\Ǆ$�      I�@�D$@Ǆ$�   !   �D���$�   �����D�\$XE���b����i����\$X���Q����X���D�L$@�v�����$�   � A         ��   ��)��2���D$P���  D���<�A���D9�tA��~�A��A�������D�a��~41�A���������A�@�����H��$�   D�P�A�   �A�D$PI���1�A�<B����L��$�   �D$D   �D$\A�@    Ǆ$�   P   ��$�   �����A�N  �������GX  ����1�����1����������+X  ����A����   Ǆ$�   !   D9d$@~�D$D����L��$�   A�@�����E����   A���]���IcPI�@H���H���@�����H9�v���t���Ǆ$�      �@���Ǆ$�      �Ǆ$�      �L$\9�$�   �<���H��$�   Ǆ$�   !   �x������xDEd$tD�d$t�����1������L��������$�   �PH��$�   ��Hc��D����ڃ���9�t
����$�   Ǆ$�   !   ����D��A������������AUATUWVSH��(�B9AH��H��|H��H�׋NE1��e]  HcVL�_H�HH��L�N�PHcGH�<�H��@ A�H��I��I��E�S�D����E��A��E�D�E�E��fD�A�A��D�f�A�A��A��H9�w��F)�H�L��L9�s;fD  E�H��I��A��A��D�A��f�A�A��E�fD�A�E��A��I9�w�E��t;St!�B�C�D�   H��H��([^_]A\A]� �C�H�u\  H�SH�HH��HcCL��   �j  H��H���N]  HcV말�������ATUWVSH�� E1�I�����D$    I�rI�ZM�Z��    1�fC�I��I���tKB�D
f��t�I�,1��D�e ����D�f�} I�,B       ��D�e D��f�E ��fC�I��I���u��   A�fA� H��H��u�H�� [^_]A\�VS����   ��~:�Z�L�YA��L�IA��L��H��D� L9�fD�@�u��1�D9�f�Au݃��ڃ�SL�Y��L�QtBfD  M��1�A� A��A��f��AH��A��A����AE�I���fA�@M9�u΃�u�1�[^�H�AE1�L�Q@ D�H��E��A��E	�E��fD�@fA��L9�u܃��r���@ A��A�ۃ����   L�I1�fY1�D  �TfA�T�H��H���u�A��1�A��f�Q�A��jE��tZH�qL�I�     �AI��1҃�	�f�A� A��A���AE�f��A��fA�� ���AE�I���fA�@�M9�u�A��u�1�f����[^��QH�AE1�L�I	�f.�     D� H��D��f��D	�E��f�P�A��L9�u�A���P���1��C���@ f.�     �A
f��f�D�A
H�AfA���fA���fD�Bt9L�BE1�H��fD�ZH��D�HI��H9�fE�H�u�E1�fD�R�f�     D�A
fA���fA���tH�BH��D  H��1�H9�f�H�u��L�I
I��I��fA�x� uM9�u���L�BE1�H��fD�JfD  H���PI��H9�fA�P�u��f�     A�   1��     F�F�E�D�fB���I����I��u��f.�     A�   E1��    B�F�D)�D)�fB���I����I��A��u���    AWAVAUATUWVSH��   �f�D$@�BH��1�L�sH��$�   1�H�D$D    L�CL���D$L    f�D$Bf�T$P��ʃ��EC       �f���f�� ���E�H���f�G�L9�u�H��$�   L�l$@H�|$0L��$�   H�kL��L�l$8I���p���t$,��)�H�t$NA��H�t$ H�t$`fD  �C������K��ȹ��  A9�r1��t$,����I��L��������   �f9��   H��H��u�1��   ���     �D�D)�)�f���H����H����u�f�oL��D  H���L9�f�P�u�1�H��H9|$ f�C�K���H�|$01�L�l$8I��fAF�I9�u�f����1�f�     A�L f�H��H��u���H�Ĉ   [^_]A\A]A^A_�D  �9���D�M�1��   ���E�D)�)�f���H����H����uܸ   �f9uH��H��u�D�������v�1����   ��f.�     �E�D)�)�f���H����H����u������    AUATUWVSH��h1��f�D$@�BH��1�H�D$D    H�q�D$L    L�if�T$PH�\$@f�D$BL�d$ �Of��D$Nf|$Pf�D$P�D$Lf�D$N�D$Jf�D$L�D$Hf�D$J�D$Ff�D$H�D$Df�D$F1�I9�f�D$DtS�H��f��t�H��M��������   1�D  �E�A�D�f���H����H��u��h����     1��f�L H��H��u���H��h[^_]A\A]Ðf.�     D�AD��f%�f=�H�A��   fE��t`E1�fD�B
f�9 L�BD�Iu9fD�JD�IfA���fA�����   H��H���P�I��H9�fA�Pu��f�fA�� �fD�J� L�IL�Y�     A�E��A���EE�f��A��fA�� �A��AE�I��D       E�fA�A�M9�u�H�A�Q����L�II��fA�8 uI��M9��5���fA�8 t�H�       ��B�  H��f�     L�QI��fA�9 �1���I��M9�u�H�       �H���    WVSH��`�A
f%�H��f=�ty�G
f%�f=�uH�W
H��H��f�x� ��   H9�u�H�\$ H�t$@H���m���H��H���b����T$ f;T$@tF�   f�< ulf�< ueH��H��u�1�H��`[^_�H�Q
H��H��f�x� u]H9�u��k��� L�L$>f���   �����D�H��A�fA9�u6H��u��f�������H��`[^_�f.�     �����H��`[^_� ����fA9�F�H��`[^_� f.�     ��t�����    1�� f.�     S�Qf���  D�AL�I1�fE����   fE��u6H�Q��D�H��fD�B�L9�u��1҃�`f�Q��   D�AfE��t�fA�� �uMH�YL�Y�E1�H��f.�     D�
H��E��fA��A��E	�E��fD�BL9�u�D�A��fA�� �t�L�Y�     fE��xML�IE1� A�E��A��f��EH��A��A��A��AE�I��E�fA�QM9�ũ���`D�A�[�1�f�� �uWL�Yf��t�L�IE1��A�E��A����EE�f��A��fA�� �A��AE�I��E�fA�Q�M9�uɃ����t��Q�H�AE1�L�Q��E��A��f��H��D	�A��f�P�L9�u��Q������m���D  f.�     AUATUWVSH��HE1�A�   D��H�ˉ�fD�d$0H�D$(    D��H�D$     fD�l$.�����)Ń�P~���  ~g��xZD��$�   E�E       ���   E1����  fD�C~iH�C��  H��f�K��     1�H��f�P�H9�u�H��H[^_]A\A]�@ ����  H�C    H�C
    H��H[^_]A\A]�f.�     ��    I�f�CH��H[^_]A\A]�D  ��$�   @��   A�   A�   A�   ��A����$�   P��A ��6  ��$�   OJ��A��uf�{ t��E1�fD�SE1�f��fD���   E���D  �Cf�������H�K1�L�S��A��A���AE�f��A��fA�� ���AE�H���f�A�I9�u΃��������H�������D��$�   ���   E�E���r�������fD  �D$,   A�   A�   A�   �����f�� ���   1�E1�1�L�\$0��    E��DD�ȉ�f�DH������H���u�����D  �CH�K1�L�k��	��A��A���AE�f��A��fA�� ���AE�H���f�A�I9�u�����fD  H�K1�L�SfD  �A��A��f��AH��A��A����AE�H���f�AI9�u��w�����uB�c�_��������    ���K�������� f�9 �At6f �f�B
f�y�H�At2H��H��H��D�@�H��fD�BH9�u��f�f�B
f�y�H�Au�H��f�8 u&H��H9�u�f�J
�1�H�    f�B�f�     H�    �B ��ÐATUWVSH��pD�I
L��E��H��fA���fA�����   D�S
E��fA���fA�����   fA���udH�Q
H��H��f�x� �c  H9�u�f�{ �S  H�CH�{f�8 �A  H��H9�u�H�    �F F       ��H��p[^_]A\�f.�     H�l$0H�|$PH���.���H��H���#����D$2�\$Rf����   H�UH��H9���   H��f�x t�H���}�����A���D$R�   H�Q
H��H��f�x� ��  H9�u������H�S
H��H��f�x� ��  H9�u�fA��������H��H��f�x� ��   H9�u�f�y ��   H�AH�yf�8 ��   H��H9�u������D  H�    �F    H��p[^_]A\��    D����H�Of��H��uH9�t�H��f�z t�H������)�H��H�������E1�H���D$(P   ���D$ @   E������$����D$Pf9D$0�4  �����f�D$PH��H���/����H��p[^_]A\� fA����4  H��H��f�x� �B���H9�u�fA����#  A��fA�����   A��E9ʺ ����    H�    E�1�f�Nf�F
f�N
�H��p[^_]A\�fA�����   H��H��f�x� u!H9�u�H��f�y� �}   H9�u��fD  fA��������H�S
�G���H�H��A�FH��p[^_]A\�@ H�H��C�F�m���H�C
H��f�{� u0H9�u��5���fD  1�f�T$P�����@ E1������     E1������     H�Q
�8���H�S
����H�Q
�9��������H��XH�I�ӋRI��fA���uH��E�SH�� 	�ux�D$D    1��$fA���twE�SD���D$D   ���  ��>@  A�� �  H��$�   D�H�D$HL�L$0L�L$DD�D$(M�؉L$ H�$� H�D$8��"  H��X�D  ��x��D$D   �ÿ���H��H�� �����	�t�D$D   1�E1���D$D   E�SG       1��q���f�     SH�� D�BA�� @  H��u�B$9B(~A��    H�uHcC$��C$���C$H�� [Ð�SV  �C$���C$H�� [�f�f.�     AVAUATUWVSH��@L�t$,��L��L�d$01�I��M��L��������n9���   ����   �F9���   �F������~WI��A�U�M��L��������~?��L��I�|�    H���K�H������H9�u���fD  H��    ������F�P����V�H��@[^_]A\A]A^��    )��F	�F�s������FH��    �����F�P����Vu��N������5���D  WVSH�� A�x9�H��L����   ����   �C9�|\���C������   �G�H�|�H���N�H���@���H9�u�C�P����S~H�ڹ    �!����C�P����S�H�� [^_�)��C	�Cu ���CH�ڹ    ������C�P����Su��u�뺉��e���@ �C������    VSH��(H��h	 H��HcRH��H��HD�H�م�x�R  I����H��H��([^����� �+S  ��f�     H��8E�X��A�@����t@H�L$,�D$,-L�QA�� E1�B�
���D	�C�
I��I��u�I�RH)������H��8�A��   tH�L$,�D$,+L�Q� A��@tH�L$,�D$, L�Q�f.�     H�L$,I���fD  UATWVSH��H��0�y�H����   �Qf��taHcFH��H��H����ɦ��L�E�H)��E�    H�\$ H���޾������   ��L�dH���K�H���^���L9�u�H��H��[^_A\]�H��.   �?����H��[^_A\]�@ �E�    �dR  H�M�A�   H�H       L�M�螲����~,�U�f�V�F�H���f.�     H��.   �����H����V���     ATUWVSH�� E����H��A�ID��L���b  A9���   D)�A�I�C9��  ���C������   ���N  �C����  �@��  �C��~�S��   ��   �~  L�c ��������  ��0   ��tH����H��� �������  �C	t�f�{  tω�����R9�u�I�غ   L���M����A�A�����C	�U���f�{  ������E����VA�������A�����~&���(�����)Ѓ�� ���Z  ��9�u�K���������N  �C��  ��  ���ɉK���������������K H�ڹ    �C����C�P����S�������H�ڹ-   �!�������H�ڹ0   �����C���C	u��u ���CH�� [^_]A\�H��������tL�C��Cf�     H�ڹ0   �������u�C�P����S~����0   ��tH����H�������C�P����S�H�� [^_]A\�)����K~d�����K������C	�����f�{  ����������� ��   ��A�I�����    ���ɉK������C����f.�     �C��u����z������q���f�{  �f��������    H�ڹ+   ������f������C�     H�ڹ0   �����C�P����S��U�����������S�J��҉K�����1����H�ڹ    �s�������������C����������C��
�C	�M���H���s��������C    ����f�VSH��hD�B�)E��HI       ��y�B   A�   �|$PH�D$PH�T$0�   L�L$LH�D$0H�D$XH�D$8H�D$HH�D$ �����D�D$LH��A�� ���tH�L$HI��H���������    H�ڹ    �����C�P����S�H���n  �H��h[^�fD  �L$HI��H������H���I  �H��h[^ÐUAUATWVSH��(H��$�   A�    �ZD�J��H��DI�A��A��   tf�z  ��  LcVIc�E9�IM�H��H����3���H)�A���L�d$ tH���   A��D�NE��M��L��A��   H��I���������tjD  I�xH��I��H��H��H�H)���0H��A�H��t?I9�t5E��t0f�~  t)H��L)�H�H��>HЃ�H)�H��uI�xA�@,D  I��뛅�~<H����L)�)҉�~,��H�LH��H��f�     H���@�0H9�u�Hc�H�|I9�u���.  E��~9H��L)�A)�E��D�V~'A���  tA��D�V���  A��   ��   �A���tZH�_�-I9�s.H���H������I9�u�F�P����V~H��    �����F�P����V�H�e�[^_A\A]]�fD  A��   t'H�_�+�D�����������A��,���f.�     A��@H���p���H��� �d����    �F�P����V�?���H��    �����F�P����V�D�N����H��� ���@ �0H�������@ D��%   =   ������V�B��҉F�������H��H�Tf�H���@�0H9�u�H�|�F��������f�WVSH�� L��I��E�H�A�gfffD��Ic�A��A��A��A��E)�A�   t#A�gfff@ D��A��A��A����D)�A��uJ       �F,���u�F,   �   D�FD9�D��I��M��WD��)�A9к����N�A�   L�҉F�����NH��F,�F�ȃ� �  ��E�F����D�OH��H��DNH�� [^_�D���@ VSH��hD�B�)E��H��xlA���|$PH�D$PH�T$0�   L�L$LH�D$0H�D$XH�D$8H�D$HH�D$ �b���D�D$LH��A�� ���t1�L$HI��H������H���
  �H��h[^�f��B   A�   뉐�L$HI��H������H����  �H��h[^ÐVSH��xD�B�)E��H���8  �  �|$`H�D$`H�T$@�   L�L$\H�D$@H�D$hH�D$HH�D$XH�D$ ����D�D$\H��A�� ����  �C%   A���|y�SA9�q����   H��D�D$<�H  D�D$<D)����C��   �L$XI��H���j�����     H�ڹ    �#����C�P����S�H����  �H��x[^�fD  ��uNH��D�D$<�G  D�D$<���C�L$XI��H���U���H���  �H��x[^�D  �B   A�   ������k���     �B   A�   ����D)S�:��� �L$XI��H������H���I  �H��x[^Ð�S������ЉC�����f.�     UAWAVAUATWVSH��(H��$�   �   �   E�XE�`��oA��I��E����    ��L�ƃ�E��AI��A��   tfA�x  ��  LcFHc�A9�IM�H��H�������1�H)�A��oH�|$ ��M�ɍ�   H����  E��A�� D  ��H��D!�D�p0��7D	�E��A��:AB�I��M�ɈC�u�H9���  E����   H��D��H)�)҉���   ��H�LH��H��f�K       H���@�0H9�u�Hc�H�\E��t	H9���  H��H)�A9���   A��o�F�����}  H9�A�����A�����s6H���H�������H9�r�E��~ A��H��    ����A�D$���H�e�[^_A\A]A^A_]�D  A��o�k����F	�a����0H���U���A)�A��o�FE��D�FtO����   A��E��~	E����   H��D�H�ZE���B0fH9�s�E�e��E�����غ����������3���E��y��   ��   ��   E�e���t<H9��#�������A������D�f�p���E��xyE�e���tH9�����������f�A��H��    ����A�D$���H9������A�����A����������0H���c����F��tkH��A���������f.�     ��   ��   t���n��������f�E�E�D��H�LH�ڐH���B�0H9�u�Mc�A��oJ�Tt��u�H��A����������f�AUATUWVSH��hL�	D�QL��H��L�L$0H�� A��D�T$8L��D�	%���D	�E������	���D	�A���  A)�D��������  fE����  f�����uf����[  f����  M��L����  D�CA����  D�CH�l$@�C���  �D$@.H�EH�p� 0D�SA�   E����   �SH��D��H)���O�1�A���  �¹gfffD�LD��A�������D)�t&A�gfff ����A��A��A����)ʉ�u�E��E9��  E)�A��   �*  D�SfD  A�����  A��   ��  A��@�2  H�ڹ0   �b����KH�ڃ� ��X�Q����C��~&�C	t ���CH�ڹ0 L         �1����C�P����S�L�l$.H9�w3�r  D  �C f��f�D$.tI�غ   L���R���f�H9��D  H�����.�  ��,t�H����������     D�Cf���?H�D$0A���x  H��x H�y��   �   H��D)���H��H���  H��   D)���H��D�CH�l$@E��E��H��A��   A�� � 1�H9�w�K��x	�J0�H��H���l  ������H9���   �SH����~���S��t���	��v�7D	���     �K�   f������`����f����    H� V	 I��1��O����H��h[^_]A\A]ÐH�ڹ0   �����C�P����S�KH�ڃ� ��P����H��H��Dc�K�  �����H��h[^_]A\A]ÿ���x����@ �׃�H�y�D�CA����������� H��D�C����������H9�wE��u	D�[E��~�.H��D�_�H��tf.�     H��D��D�_�H��u�1������f�     H������������ H9�������m���f�H�ڹ-   �����/����C��������f�H�ڹ+   ���������������fD  A��D�S�     H�ڹ    �S����C�P����S�D�C����H�ڹ    �0�������A��   H������������H�JT	 �� �  I�������>���f�f.�     AWAVAUATUWVSH��   H�-&T	 L��$  A��H��D��L��A�� `  ��?  1�1ҋ f��$�   �H�|$pD�d$xǄ$�   �����D$8H������H�D$|f��$�   Ǆ$�       Ǆ$�       ��$�   ��$�   H�s��t��%t7H�T$p�=M       ����KH��H�s��u⋄$�   H�Ĩ   [^_]A\A]A^A_� �CL�l$pH��E1�H�\$`D�d$xE1�H�D$|����M�]H�\$(H�_�Ȅ�A���0  �P���Z��  ��HcT� H����    I�I�wA��A���  L��I���������4����     A�I�wA��Ǆ$�   ����A����  H�L$`M��D$`I���   �����D  E���'  �L$x@�GH���D���fD  �D$xI��I�W��� ��D$x��  �*L��H�L$@�|$@������]���E����  �L$x   �G�fD  �G<6��  <3�6  A�   A�   뀃L$xA�   �G�l���f.�     I�wI�?H��Q	 H��HD���$�   ���  Hc�H���;  M���H������I������I�wA����  A��A�tA����  A��u��H�L$`A��ut[H��M��D�������I���q�����L$x�   I�wA���,  A��IctA����  A��uH��H�L$`H��H��?H�D$hL��I���Q��������D$xI��I�W��� ��D$x��  �*L��H�L$@�|$@���������f�     �D$xI��I�W��� ��D$x��  �*L��H�L$@�|$@���������GA�   A�   <l�����H�_�GA�   �����f��GA�   A�   <h�����H�_�GA�   ����D  �GA�   A�   �����D$xI��I�W��� ��D$x��  �*L��H�L$@�|$@���������     I�I��A��Hc�$�   ��  A���  A��t
A���.  ������fD  �L$8�: N        L��H���|��������    E��uD9d$x��  I�I�wM��x   H�D$h    I��H�T$`�����f���fD  L��%   ������N���Ǆ$�   ����I�wA�H�L$`M��   I��f�D$`���������D$xI��I�W���D���H�T$(H�L$@�D$(L���|$@����������f.�     �D$xI��I�W���W���H�T$(H�L$@�D$(L���|$@���������D$xI��I�W���y���H�T$(H�L$@�D$(L���|$@�����z���f.�     E����   �L$x   �G����fD  E���  �L$x   �G����fD  �D$xI��I�W������H�T$(H�L$@�D$(L���|$@���������A����  �GA�   �F���@ M��t�A��������   A�I�W��A��"  �GI��E1�����E��u(�L$x   �G������    E���s  �    �G������    ��0<	��   A����   E��u-A�   M��t�A�����   ��A�DA�A��A����   A���   DD���f.�     H���D����GE1�A�   �X����2�r  H��A�   A�   A�3   H������H���6  �����f�����Ǆ$�      D�����D$x����H�����L��%   H����������A��0�GE�������GM�]A�   Ǆ$�       ������M����4u�H�_�GA�   A�   ����I�H�L$`�����I�H�L$`�����L$x   D�T$<L�\$0�D$`    ��6  L�L$(H�L$^A�   H�P�����L�\$0��D�T$<~�T$^f��$�   �O       �$�   �5�����H�L$`����H��H�L$`�b���E��u4�L$x   I��E1��\$|�G�����H�_�GA�   A�   �����Ǆ$�   ���������SH�� 1ۃ�~�   ����P9�|���'  �H��H�� [�WVSH�� A��H��H��~m�   1�fD  ����HA9����l'  L�F�D�H��H�@E��D�IH��tI��E�H�H��E��D�	u�H��tH�H�� [^_�f.�     1��f�f.�     �   H�ȋI���HH�H��P��'  @ AWAVAUATUWVSH��81��r9qI��I���g  H�Z��1�L�iHc�H��H�<+L��H�E ���A�ƉD$,��   ��I��M��1�E1�I��A�K�I��E�B�H��H�H�ȉ�I)�H�� M)�M��E�B�I�� A��L9�sƋE ��uCH�E�I9�s5D�]�E��u,H��L)�H��H���H��H�T��D�E��uH����H9�u�A�t$L��L����+  ����   A�FL��1҉D$,�    H���H��D�C�L)�H)�H�A�H�� ��H9�s�Hc�I�T� D�
E��uAH�B�I9�s3D�B�E��u*H��L)�H��H���H��H�T
�����uH����H9�u�A�t$�D$,H��8[^_]A\A]A^A_Ð���AWAVAUATUWVSH��   )�$�   A�9��H�͉�$�   L�Ã��M��A��������4  H��I	 Hc�H����11Ƀ� ~�    ���9����$  H��I�ƍF�M�F��H�L��L���    �
H��H��I9҉H�s�L)�H����H�I�D���H��E��D����  �D�j���t�Mc�A�V��C�D�A�Ճ�A)�L���  D��$�   ����$�   ��  E�P       ~E����   L���5%  H��$   A�   H��$(  H��H	 �    �m���I��(�$�   L��H�Ĩ   [^_]A\A]A^A_�H��$   A�   H��$(  H��H	 �  ����#���I���H��$   A�   H��$(  H�qH	 �  ��������I��뇐H��$�   L��D�L$,�++  D�L$,fI~��qH	 L��E��H�� G�)���� A�@���  �?H��H�� I	׺   fIn��\'H	 D)��Y$H	 ��IЁ�5  ���X�f���*��YH	 �X�~f���*��YH	 �X��,�f��f.�T$,��  ��E���D$\   ���H�� I	�M��L�|$pM��D�|$,A��w/H�}W	 Ic�fIn���f.��V  A���D$\    D�|$,D���D$H    )��ʃ��T$@y�   �D$@    )ʉT$H�L$,���N  L$@�L$d�D$0    ��$  	��  ��$  ��  �  =�  A����$  �
  �   ��$  �D$`   �   ��$  �\  �D$,�$  �H�D$|���L$8��A!�����
  ��$�   L�T$hD�D$xD�L$P����D�L$PI�ǋED�D$xL�T$h���D$Xt!�L$X�   ��I����   )ȃ�D��D$XE���A  �D$,D$X�D$P�/  Ǆ$�       D�T$\�T$pE��t�4F	 f.��@  f(��X��X2F	 fH~�fH~�H�� ����  @H�� H	ЋT$8���J
  D�\$8f(�E1ҋ|$`fHn�H��U	 A�C�H����,��"  ��E	 I�Ǆ$�       �,��^͍B0A��\�f���*��\�f.���   �-{E	 f(Q       ��\�f.��  ��$�   ��D9؉�$�   ��	  �OE	 �,f(��\�f.���  ��$�   ��D9؉�$�   ��	  �Y�f��H���Y��,��*���0�G��\�f.�v�f.�A�Zz�Q  �D$P   �D  A�F    �6�����L����  ��$�   D��$�   A)�A��1���Ǆ$      f���*�L�T$P�Y{D	 D�L$8�,ȃ���$�   �s���D�L$8I�ǋEL�T$P���D$X�  ������D$`   Ǆ$      �D$|�D$8fD  E���  �D$,9E�
  D��$  H�H��S	 H��E������  �D$8����  ����  �Y�C	 fIn�f.���  H�D$0    ��1�I�A�1�D$P    H�L$0�u  H��tH���h  L���`  H��$   � H��$(   �tH��$(  H�8�D$PA	$�&����D$\    ���� ��$  E1����������E1��D$`   �D$|�D$8Ǆ$      �}����     �L$`���d  �UD)�D�ɍF)�$�   9��7  ��$  �N�����$  D��)Ѓ����t$8����$�   ����t9��  �t$H�|$0D$@��t$P�D$H�   �z  H�ƋL$P��~&�T$@��~9щ�N�)D$H)�)�$�   �L$P�T$@�D$0��t1�T$`����  )���A����  L��D���}   I��f.�     �   �  A���T$dH��H�D$0����$  A��A!Ņ��_  E���h  �   +l$@�T$H����ꉬ$�   ���~L���!  I�Ƌ�$�   �T$@�~H�L$0�k!  H�D$0��$  �D$\@R       �ǅ��.  D�\$8E���   @���  D�T$8E���"  ��$  L���D$P   ������f���*�f.�z�)����l$,����f��L$,�D$d    )L$H�ىL$0����D  ��$  �D$`    �J���D��$  �   E��O�$  ��$  ��$  ����$�   ��A!��L$|�L$8������    �D$H1��|$0�D$P������  E��H�D$0�  �D$d    H�|$0�G�D$x��H��l����v���@ D�L$`E���R  �T$P��~H���    H��D�D$dH�t$@E����  L��$  L�d$@Ǆ$�      L�|$HH��$   ��   L���  ���$  uH��$   � �D$@��T$X��	  E���<  D�$  uH��$   � �!  I���~�|$X�  @�o��D$89�$�   �;  E1�L��
   �  E1�L9�
   I��H����   �  L��E1��
   H���u  I�ă�$�   I��H�\$0L��H�������H��L��h0����  H��L��   A���   �HI���������H��L��H�D$@�  L�D$@�������f.�     ��  H��I��� ��$  ������t$0�D$8����)�9�}��+T$01��D$0T$d�D$8����  �t$H��$�   D$@��t$P�D$H�����D  H�T$0L���  ��������l$,E1�L��
   �f  D�l$|I��E����!ǋD$`����  �D$|@���D$8�����f�     Ǆ$�      L���\$8L�l$0�"�    L��E1��
   �   ��$�   I��L��L������H���h0@�o�9�$�   |�E1�\$S       X����  ��A�F�W���  ���  L9���  �P�H��H�G���9t���D$P    �H�L$0�  �\$,��H�������M�������I9��z���L����  �m����D$`    ����fIn�fInL$,Ǆ$�      �^�I������,�f���*ʍB0A��Y��\�f.�ztt��$�   D�D$8D9���  ��<	 �f�     ��$�   D9��`  �YÃ�H����$�   f(��^��,�f���*ʍB0�G��Y��\�f.�z�u��D$P    ����H�L$0E1��   �e  L��H��H�D$0��  ��������\$,���B���H�D$0    1�����Ǆ$�      �   ����f(��X��X�;	 fH~�fH~�H�� ����  @H�� H	�f(��\�;	 fHn�f.���   fW�;	 f.�w�fI~��D$X    �D����T$0L���  I���@�����H��D$0�  L��H��H���d  L��H���	  D�D$0I��E����������� �D$X����  ���D$P   �k����G��L9��h  �B�H��H�W�<9t���D$P    ��;����D$,A�1�D$P    �w���H�D$0    �   1�������Y�L��1���:	 Ǆ$�      f(��fD  �Y˃�D����$�   �,���tf���*�D���\�H����0�G���$�   D9�u��:  �b:	 f(��X�f.���  �\�f.������f.�z��  �D$P   A�J��     H�ǀ�0H�G�t���D���L��   �  H�T$0H��I���  �W��� �V���u	���K���A�F���D$P   T       �  ��W�H��H�G���0t��5����T$XL�d$@L�|$8L��$  �|$\L�|$H���b  A�~��  �|$X��  H�\$0L��$  L�l$@H�|$8�FE1�L��A�l$��
   �P  L9�L��
   HD�E1�H���6  H��I��H��I��L��������h0L�gL��H���  �����9H�|$8L��L��L�l$@L��$  �  ���D$P    H��H�D$8I��@�(H�t$@�B���Ǆ$�       �D$H+D$8�D$P�����A�Z�v����E��9�$�   ������D$d�D$d   �D$H�D$@��������J����N��  H�VH�HH��HcFL��   �	!  �   H����  H�D$@������L$8���
���D�\$|E���R�����7	 A�������7	 �Y��Y�f(��X�7	 fH~�fH~�H�� ����  @H�� H	�����A�0���G�L��������9L�d$@L��$  L�|$8L�|$H��   H�D$8��I���D$P    H�t$@@�(�����L��I��L�|$HL��$  H�������X��G�f.�����zu	�������D$P   ��������   H�D$8�D$P   A�~H�X�.���A�~ �D$XED$P�D$P����A�F���O����D$P    ����H�D$8H�xH�D$8I���9   H�t$@� 9�����E��9�$�   �������� L��   �#  H�T$0H��I���  �� ��   ��9t��l$\�D$X    ��1�7���E1�H��
   �Q  @��H�ƋD$|�D$8���������A�~��Ѓ��D$P�Z���L����9�|$\L�d$@H�xL��$  L�|$8L�|$H�T$P����E��~}�l$\�D$P    ��1U       �����A�~ �G������(���H�D$8�D$P    H�X������D$P    A�J�t���H�D$8�D$P   H�X����u
@�������D$X    �H���A�~~�D$P   ����A�~ �   DD$P�k���E1������f(������������AWAVAUATUWVSH��8I��H��L��$�   M����  H�5�C	 L�0�~0 ��  I�E I�$    �H��0�-  H��E1�fD  H��H���H�A����0t���E��< ��  E����  D8���  H�BM�N�H��I��A8���  E��E��u�������#  ��0H��uH�����0t����E1҄�H��A�   A���3  A8�A�   H���C  H��D��D$$    t	)����D$$A��P�x  A��p�n  E��I�] �  H��1�H)�����~ ��������Q  A�~ I��H�@H�D$(�a  A�   �f�I��C�| I�Au�H9��G  K�E1�L�t$(E1��&�    D��A���L������A	�H9��   �C�L�{�:M�F��  A�� u�I�NE�A�   M���C�I��E1�1��f�     A��H��E1�1��f�H��D�JH�ZB�< u�E8������H����  D������f�1ۉ�H��8[^_]A\A]A^A_�H�Ѐ�PH��H��t��ptA�   �D$$    E1�1��K �D$$    A�   �C<+��  <-A�   ��  �CH�SD�1�H��E�Y�A����  H�W�E��HD�E��I�E �`������E���E���E�|  ����  ����  ���1  �] �ރ����������1ɉ���V       tfD  ����u��d  ��I�$�x~�N�H�PH�L������H��H9�u�A��9�~A�    Ic�D��)�A��D�D��E�   H��$�   �����f.�     �  �p���fD  L��L)�H9�� ���A�Ã�L+D$(E��u I��E�EA��A)�A9���   �    ��  �D$$9E�7  �E�L$$9���  ��)�9���  �U���b  ���<  ���  L���^  �  �P   � "   �����f�     H�SE1��D���@ ���8  ��u�D��$�   E��t�1��  I��H�      I�E�EH��$�   M�,$�b   ��2  � "   �y����    ������f�     D��L��)���  ����t0�K�H�T$(A�   �   ��A����H�D��t���a  �   ��L����  \$$����L���`  �  ��   � "   �����E1��K��� H�PE1������@ H�BA���R�!f�A��   ��   E�H��C��E�LS��D�D�ڃ���v�D����E��DE�DL$$�����   ��t!�E���+  ���5  ���6  ��H��$�   M�,$�t$$�0�<���f.�     A�F����  I�NH��8Ct�  �H��H��E8���  D�	H��D�E��u�A��H�À< �����H����< I��u�����f�     ��L��D)É��  )\$$I��H�@H�D$(�P���D�s���tE�   L�|$(D��D��   �����H���A����E�L��)��  �E�   �D$$�����E��t�D��L����  ��문   +�$�   ��$�   ��$�   �W       ������L��Ic}荊����I��H�@�Z  A9}��t2�D���    )��9�~�   L���  �D$$�D$$9E������!   �e�����$�   �������H�|$(A�E   �   �����D��$�   E������������E1�����M�EL�t$(�    E1������D��$�   E���J�������D��$�   E���4��������D��D$$    �����@�������H�D$(8�����������9���������G����V�L���  ��������E�,�����$�   �������������L���u  ��������   �����U �"   ��9��?�����A�   ����1�A��Hc�D���Ã�!�����D$$    �+���H�BD�[�b����ATUWVSH�yI��HcI����9���   H���H��L��H����   D�L�CA�    ��A)�A��M9�v7H��A� D��H��I������D	ЉF�E�P�A��M9�w�I)�I�C�H��H�|�E��D�tH��H)�H���JfD  A�A    A�A    [^_]A\�f�     I9�H��v��     �I9�w�H��J�H���x��A�yt�[^_]A\� f.�     HcAH�QL��L9�s/�I1���t�@ �
��uH���� I9�w�������    1�Ð�������������   �0   H��� L��*	 �     D�BH��D�A���u�   �a   L��*	 f.�     D�BH��D�A���u�   �A   L�Y*	 f.�     D�BH��D�A���u�Ð���������AWAVAUATUWVSH��HL�5�8	 A�~0 H��$�   ��  �������Hc҉X       D$<H��$�   M�,�I�ULE�L�I�]�A�E�    �I��A�B����v��0�T  A�RE1�E1�1�L�l$0��H��H��I�B��   ��A�����   �� �H  D9���   H9�sUA��OA�   �A�    H�D$(E)�I��A��E)�@ E�aD��I��D����D��	�A�Q�D����A�L9�w�H�D$(L9�A�   wz�PI��I�B���g�����L�l$0�   ��   H��H[^_]A\A]A^A_�@ A����A�������	щ�D  L9�v��F�    1�H��A�   ��fD  H�n��F�    A��E1�H��A�R�� wf�H���P�� v��0�P����P��߀�X�@����x �6���H���-����    ��)L�l$0�R  ���J  H��$�   I��L�H9�sKA��E�A�   �    E)�I��A��D)߉�@ E�Q��I��D����D��	�D����A�A�A�L9�w�L9���   L�ǥH9�s�f�     H���G�    H9�s�A�E���t�vfD  H�����ufI9�u��   �   �|����A�B���<X�����A�R�� �����I������f�     L�D$0H�T$(�Q���L�D$0H�T$(����f��   �!���fD  �|$<A�E����d����    �����)���!�A�E��K����    I�B��)tA�R��u	����tH����)u�H��$�   H��   �����������VSH��(�D� ��Hc�t8��tX��uH�� �   �Ӌ� ��t��tH��([^���    H��H�	� H��H��([^H�%�� �     �   �Ճ ��t��t��ƃ ��t��Y       �H�ȃ H�� ��H��� ��H�   蚵�����    �@ f.�     SH�� �   �p� ��tH�� [�D  H�� H�b� ��H��� H��H�� [H��@ f.�     VSH��8��1��������	<H�ł Hc�H��H��tyL� �=�� L��uUH�D$(H��� �3� H�D$(�<��   ��C�H�H��'   H�����   H!���  H��t�=�� �p�Xt�H�@    H��8[^�D  H�I� ��   ��S�H�&y Hc�H��'   I��I)�H��L�ɉ�H��H�H��   �h���H��H��� 눐f.�     SH�� H��H��t,�y	-1������HcSH��� �=� H��H��H�tH�� [ÐH�� [�F  fD  H�� H�� [H�%�  f.�     UWVSH��(�qH��Ic�Hc�L�I1�fD  A��H��H�H��A��H��H�� 9��H��H��t9w~%Hcƃ�H���\��wH��H��([^_]�f�     �G�H����H��H��t�H�HHcGH�WL��   �$  H��H���������    SH�� �˹   �����H��t
�X�@   H�� [�f.�     AVAUATUWVSH�� HcyLcjH��I��D9�}��H��Ic�I��Lc�B�/1�9]��M�m���H����   H�pHc�L�$�L9�sH���    H��I9�w�I�VH��N�,�H�|� L9�r�bf�     H��I9�vPH���J���t�I��I��E1���M��I��E�A�E�2L��M�M�rM�M��E�F�I�� L9�w�H��I9�E�Zw���~"E�D$�I�T$�E��t�f�H���
��u��u�XH�� [^Z       _]A\A]A^�D  f.�     ATUWVSH�� ��H�ΉӃ���   ��H����tRH�=v H����   L�%� H�����t2H�7H��t8H����t�H��H���q���H��H��tlH��H��������u�H��H�� [^_]A\ù   �����H�7H��tM�= u�L���T� �fD  H�i!	 ��E1�H����)���H��H���G���1�H��H�� [^_]A\�H��H�������H��H��H�t�H�     딹   �T���H�=-u H��t�=�~ ����H��~ �ʐ ������   �?���H��H��tH�   q  H�=�t H�GH�    �H��t     1�������    AVAUATUWVSH�� H�͉�A�֋ID�m���EA�A�]9�~f����9�������H��I����   H�x��~#�V�I��H�D� A�     I��I9�u�H�|�HcEH�uA��H��tiA�    E1�E)��L�ϋL�OD��H�����D	�A�I�D�F�D��A��H9�w�A��E��D�GAE݃�H��A�\$�"���L��H�� [^_]A\A]A^åH9�vإH9�w���f�LcB�AD)�u1N��    H��N�	J�T
�L9�sH��I��D�E9t�����f�UWVSH��(HcB�YH��H��)��  H�QH��    H�
H�L�	H9��  H��H���998t���   �N�g���H����   HcVH�N�XE1�L�]L�PH�<�H��HcUI�,��
�    L��L�II��A�s�I��A�Q�H)�L)�I�Љ�A�R�I�� A��L9�w�L9�v=M��D  I��A�Q�I��L)�I�Љ�A�S�I�� A��L9�w�H)�H�W�H��M�T�I����u I��A�����t�X[       H��([^_]�fD  �    ����H��   H��H������f�1��i���H��t�H�@   H��([^_]� SHcAL�Y�    M����E�J�I�Z�E��A��D)�A��
�A�   D��1�D)���  �?H�� I9�sA�R���A�HA��A	�L	�fHn�[�f.�     A��I9�s[E��A�R�tY��D��D��D)���A�щ�  �?A��D��D	���I�J�H�� I9�sE�B��A��D	�H�    ����H!�H	�fHn�[�1�E��uD��  �?H�� H	�fHn�[�D��D��1���  �?H�� �f.�     WVSH�� �   fH~�H��L���$���H����   H��I��H�� A����A���� ��E��A��   ���  EEȅ�tjD��E����   �    E��D)�A��D��A��A��E	�D�PE1�E��D�HA��A����D�@tEB��������5   D)ډH�� [^_�f�     A���@   A�   D�Y A���D�Hu�Ic�A��A��2  �T�D���A)�D�H�� [^_�f�     �X�i����     H��H�J��҈tH���Q�H���҈u�Ð������������AVAUATUWVSH�� H�Ήպ9��8A�HD��D�ˉ�������)ʃ���   �   1� ���9��������	Lc�$�   �X�@   ~{H�^	D�m�N�t.
H��H��D�F��
   H��A��0�����L9�u�K�T,H�9�~/��)�H�t;fD  H��D�C��
   H��A��0����H9�u�H�� [^_]A\A]A^�f�J�\&	�	   �@ 1��R���f�     UWVSH��8H��H��H�T$(����H�T$,H��fH~�fH~��q����G+EfH~�fH~���D$(+D\       $,��~2H������H�� �H�� H	�fHn�fHn��^�H��8[^_]�D  fH~�����H�� )�H�� H	����    L��A� D�X�D�P A��AB�D9�u"H��D�J�I��E��uո   L���    1�� f.�     WVIc@I�p��H����Hc�H9�H�T�s*H�ϥH9�w�L)�H��H��H�L�H9�v�H���A�    H9�w�^_� f.�     HcAL�IA��A��D9�}>M��M9�ssA�@�I�P���uWH��L)�H��H��H���L���H��D�E��u4H9�u��Ic�D9�M��~���t�E���D�������¸   A9�t��@ �   �f.�     1�Ð������������H��I��t�9 u���9 tH��H��L)�H9�r��1�Ð�������1�H��tf�9 u
��f�<A t	H��H9�u�Ð���������������%Ƌ ���%�� ���%�� ���%�� ���%�� ���%v� ���%f� ���%V� ���%F� ���%6� ���%&� ���%� ���%� ���%�� ���%� ���%֊ ���%Ɗ ���%�� ���%�� ���%�� ���%�� ���%v� ���%f� ���%V� ���%>� ���%.� ���%� ���%� ���%�� ���%� ���%։ ���%Ɖ ���%�� ���%�� ���%�� ���%�� ���%v� ���%f� ���%V� ���%F� ���%6� ���%&� ���%� ���%� ���%�� ���%� ���%ֈ ���%ƈ ���%�� ���%�� ���%�� ���%�� ���%n� ���%N� ���%>� ���%.� ���%� ���%� ���%�� ���%� ���%և ���%Ƈ ��]       �%�� ���%�� ���%�� ���%n� ���%^� ���%F� ���%&� ���%� ���%� ���%�� ��SH�� ���T   ��H�IH��H�H�� [ÐH��s ��     H��H��s Ð����H��$	 H� Ð����H��$	 H� Ð�����%�� ���     UWVSH��(L�ˉ�H��L��L���Є HcHc�H��H�H=���P�+��xH���,� 1�H��([^_]�D  ��H��9�O�E1��1� ��u����+H����� �   ��@ H���� �"   H��([^_]�f�     SH�� H�҉�tH��r ��r H�� [ÐH�=�r  u�   �� ��r H��r H�� [��     UWVSH��H��r ��H��H��t:H�H��t@�h�8�� L�H�t$0H��	 H�or A���l$(�|$ �_����H��H[^_]�D  ��� L�H�t$ H��	 H�4r A���,����H��H[^_]�f�H��t1��    �f��   �f.�     H��t1��    �f��   �f.�     H��tH��t��1�ø   �f�     H��tH��t	1��    ø   ��    H��t��u1��@ �   �f.�     ATUWVSH�� �   ��M��w`��L��uc�  H�ý�� �f�H)�t*H���� H��HB��8  ��H���^.  �)  H)�H9�w�1�M��tI�$    I�D$    H�� [^_]A\��y  H���@ H��t��w���    �(   t1�� �   �f.�     WVSH�� H��H���  H��t	�:�  ��   �   �����H�ø   H����   �����1�1�H�=�� E1�A���^       �H�H�C    �C    ��1�E1�1�H���   A������H���   H���   H��tVH��tDH�=с H�K��H�Kp��H�K@���Ch    1�ǃ�      �����H�H�� [^_��    ��� H���   H��t	H���� H�������   H�    H�� [^_�f�     �   H�� [^_� �(   H�� [^_� VSH��(H��H� � �{  H��t61�H�;�tH�� �  ��H��([^�f�     1�H���v�������f��   ��f�     UWVSH��8��H�Ή�D����   H�L$ �-(  H��H�D$(��   H�5�� H�|$ E1�A��H���   �փ��*  �    rG=�   �
  =  �=  ��   1�H�L$ �_� ����  ������t�T)  ����   ��H��8[^_]ÐD��H�=*� ��=�   ��   =  ��   ����Ӄ���H��8[^_]�f�     ���H�=� tq����   �   H����=�   �  =  ��   ����   ��t	�(  ��ue�   �������V������N�����)  �D����(  ���3  �(   H����=�   ��   =  t�1ۅ������X(  ���   �   ��H��8[^_]Ã��   ���������   1�H��    �ׅ�E݉�H��8[^_]É�H����=�   tS=  t���=���1��;�������   1�H���ׅ�u1������   ��   �������t�'  ���^����   �����@ �'  ��uG1�H��1��ׅ��É�H��8[^_]û   �����@ H�L$(��~ ��u�(  ����fD  ��������r(  �_          ������3'  ���7��������fD  AWAVAUATUWVSH��8L�%�} H��$�   I��A��D�D$,L��L��A����+H�-�} 1�D�+H����E��D�D$,x��H��8[^_]A\A]A^A_�D��L�������H���A�ԅ�uH�����������    AUATUWVSH��8H��H��t~H�H��tvH���t>H���   H�kp1�A�����L���   I��L�d$ �'�������tq��H��8[^_]A\A]�f�H�� �   �_  H�>�t9H�Ҙ �  ��H��8[^_]A\A]ÿ   ��H��8[^_]A\A]�f.�     H�    1��D  L�kL����} ����   �C9C~3H���   M��I��   �,���L����Ǹ   D���| �A���f�H�    M��I��   H���   �����H���   H�5�{ ��H���   ��L���<| H�5�{ L����H����H�K@��H���1��������H���   M��I��   �   ���������f.�     VSH��HH��t%H�H��tH���tz�;�����   tH��H[^� �   H��H[^�@ H�sH���{ �C��tL�S����   �����S�CH���x{ H���   L�Kh�   L�C@H��H[^�����1�H��H[^�@ �C9C~XH���   L�Kp�   A�����H���   H�D$ ������u=�S�C��t	)��C    ���C   �C�s����     H����z 1������D$<H����z �D$<� ���f.�     WVSH��@H��t$H�H��tH���tw�;�����   tH��@[^_Ð�   H��@[^_� H�sH����y �C��tL�{����   ��C    �CH���Hz H���`          L�Kh��L�C@H��@[^_����1�H��@[^_�D  �C9C~MH���   L�Kp�   A�����H���   H�D$ �������u2�C�{��t	)��C    �C    �{�v���H����y 1��"����D$<H����y �D$<����D  ATUWVSH�ĀH��H��H��t[H�H��tSH����  �;�����   u/H���   H�sp1�A�����H���   I��H�l$ �%������D$<tH��[^_]A\�f��   H��[^_]A\�L�cL����x L��C�y H���   I��I��   �������D$<u�H�D$<H�\$@H�D$PH��   H�D$`H�D$@H�|$HH�D$h�x   H� H�D$p���h   H�T$`H��H�����  ���D$<t=�H   H�T$pH�H�L$h�T$`�D$<�1�������������D$<����H������f�H���   H�ChA�����1�H�D$ L�K@�����D$<�f�     AUATUWVSH��HH�H�kH��H���}w �{��tZ�G�H��C��w ��u H���   L�Cp�   L���   �Z�����uH�N�]  ��tH�V�H��H[^_]A\A]�fD  �C=���?t&���CH����w H�N�  ��u����     H���   H�{p�C���?A�����L���   I���   L�d$ ������A��uI�CM��I���   )CH���   ������u�C    �{����D$<H����v H�V�D$<��<���H����v H�FD�(�'���f.�     ATUWVSH��   H��H��H���4  H�H���(  H����P  �;�����   ��   E��L���  ��  �����H9��  ��H���   H�kp1�A�����L���   I�a       �L�d$ �%������D$L��   �CM��I��   H���   �������D$Lu~H�D$LH�\$PH�D$`H�����H�D$pH�D$PH�|$XH�D$x�  H� H��$�   ���  H�T$pH��H����  ���D$L��   �p  H��$�   H�H�L$x�T$p�D$LH�Đ   [^_]A\�f.�     �   H�Đ   [^_]A\��  �����H9Љ����������������D�L$<L�D$0�����������D$Lu�H�L�D$0D�L$<����f�H���   H�ChA��1�H�D$ L�K@������D$L�D���f�     E1������     A�   ���������H��8H�L$(��t �T$,H� ��*!Nb��D$(H�� H�H�KY�8��m4H�H��H��H��H��H��8�f�     ���CLi�  �I��������)�Hc�L��@ f.�     SH��0���CLi�  �I��������)�H�L$(Hc�L���s �T$,H� ��*!Nb��D$(H�� H�H�KY�8��m4H�H��H��H��H��H)�H9ں    HG�H��0[Ð������VSH��(H�ι   H������H��H��t=H����     �   t	1�H������AH��H�A    �A    �A�����H�u
H��H��([^��v���H���UWVSH��(H�H�CH��v+�   ���;��u>�S��u1�H��([^_]���r �C��H���H���H�ø   H��u�H��([^_]�f��C��uIH�{ trH�=�s �   ����������t�H�K���ׅ�t�=  �   ��   E��f�     �k�Cr 9�u�����;�$   �{�Y����C1��N��� 1�E1�E1�1���q H��H��t1��H�K�h����b       �q �]�����q �   ���   E������@ ATUWVSH�� �����H��H��t&H��1�����H���7���H9�vH)þ����H9�HF�H�H�CH��v6�   ���+��uL�S��u1�H�� [^_]A\�D  �Vq �C��D  H��H�������H�ø   H��u�H�� [^_]A\ËC��uFH�{ toH�-lr �   �����t�H�K���Յ�t�=  �   ��   E��x����     D�c��p A9�u�����+�$   �{�L����C1��A����1�E1�E1�1��\p H��H��t1��H�K�k����8p �`�����p �   ���   E������@ SH��0H�H�BH��vD�BE��u51ɇ
1���tjH��0[�@ ����H�¸   H��u�H��0[��     �
�   ��tˋZH�T$(��o H�T$(���   9�u��B��u$�B������    H�J��p ������낃��B1��u���D  f.�     VSH��(H�H�CH��v11��   ��uB�C1���u	��H��([^��do �C��H��([^�H�ھ   �����H��H��u���H��([^Ã{t�   뺋s�$o 9�u�C1��f�f.�     H��t.��(   ��u!��H��������t1�����H�D �H�1��H��������@ VSH��(H�H�CH��H��vH�KH��t�_n H������H�    1�H��([^� 1��    ��    H������fD  H��tH��t
����1�ø   �fD  �   H��t��w����	�1���D  H��tH��t������1��f�     �   �f.�     c       H��t��w���(   �    E!��f��   �f.�     ����1��fD  �   A��A��A��u����	�1���f�����1��fD  ������1��Ð1�H������fD  1�� f.�     1�H��H�H��t1���H�H��t���@ 1�H�H���������@ f.�     1�H�����Ð�����1�H�H��t1��:�m@������     WVSH�� H��H�� �z���H�5�[ H��tnH;>u�G�    H9;H��t;H�^H��u�    �   �`���H�8H���@   H�FH�K1��t����	f�H��CH��� �M���H��H�� [^_�f��    �   ����H��H�8�@   H��Z 묐f.�     H��(�:m ����e� tH��(�������L��Z M��tFI��L��Z t<I��E1��L9�t+L�@�M9�r"K�H��H��H��L�H9Jtw�L�HM9�s�1��I;Ju�I�ÐH��f�f.�     ATUWVSH�� H��H���  H�=[Z H�LZ L�%UZ H9���   H�-Z I�       @H��L��H�Z t4H�Z    �   H���#���H��tH��Y H��L��H��Y u�H��t���H��t=H��H��H���I;\���   H��H��u�L��I���   L�I��H�������I��H��H��I�\$I�,$H�=�Y H�� [^_]A\�H��u9�   �����H��I��tH�ZY    H�cY ����1�H��H�� [^_]A\�H�GY H�XH��H���?���H��I��t�H�Y H�!Y �����I�4H9�uI���]���I��I)�H��H��H���5���D  WVSH�� Hd       ��H�7� �����L���  M��unH�KPH��t�P���H�KXH��t�B���H�K`H��t�4���1��<   H���H�H��X H��t~H���  H��X H�΅ H�� [^_�*���f.�     L�QX M��t�I�x�H�5IX 1�H���f�H9��i���H�H�H9��\���H�
H��I��I��N;Ttr�H�P��H�X H�X �H��I9�w4H��H�=�W ����H���l���H��W     H��W     ������H��I)�H��I��H�H�L�������f�VSH��(H��H��� �K���H�TW H����   H9�u	�   �H��H�CH����H9���u�H��tD�ntH��� H��([^�<���H�N����H��H�FtH�CH��������H��V �� �   �� H�.� I��H������룐H��1��f�     SH�� H��H�I����H��tH��H�� [����H�� [��    SH�� H��� ����H��V H��tSH������H��H���  t3H���  H��H�~V t\Hǃ�      H��� ����H��H�� [�1����     ��  �   ����H��H��t�H������H��tH���  � H�V     � H��1������@ WVSH��   H��H��t������tH�����H�Đ   [^_�H�|$ 1��
   H�5�� �H�|$H�C   �H�\$ ��f H�S'A�
   ��� i �|$G t2�(   �fD  H��H��kt�< ��u��juH����f �3����'   Hc��D 
�BH��D  ��f�WVSH�� H�BU �M���H�pH��H���.����=(U ��u4������U    H���e       ���H��tH���@���1�H�� [^_�fD  ��tֹ   ��� L��T A��H�b� H���W����D  UWVSH��H�=�T t�Z����� ��f H��H��tH��H��H[^_]�f.�     ����H�=À  H��t�H��t��@D   �Xe E1�E1��   1ɉFp�e H�NhH�F8����H�F0�!���H�e ǆ�       H�F(    ��H���e H�����D$0   I��H���D$(    L�N(H���D$     ��d ��tIH�N(�e H��� ǆ�       ���   �F@��σ��F@��e ��tH��H��H��H[^_]��S����f.�     SH�� H��H��t3H��� �g���H���O���H��� H�������H��H�� [��    1�H��H�� [�D  AWAVAUATUWVSH��(����H��H����   L�`hA�   H�->� L�������GH����   E1�1��@ ��;_HsqH�GX�ހ<0 t�H�GPH��L�<��"  H�UR H�<�H�GPH��    H�GX�0 v#L��A�   �l���H�%R L����L������H�����$  ;_Hr�L���?���E��t
A���R���H��([^_]A\A]A^A_�L��H��([^_]A\A]A^A_�����    WVSH�� ��uM����   �   H�� [^_Ã���   ��u�3 ���t���c H��H��t��@@0��   H���  H����  H�K(H��t$H�5bb ��H�K0H��t��H�C0    H�C(    H�K8����H�Kh�o���H���   ��   H���Y�����   @ H�Q H���D�����b H��P     �.���f.�     H�����   ��a H��Pf        ����f�H�H0���   ����   H��t��a H���  H�C0    ǃ�      H����   �CDH�{8H�sh��   H�K(�ﾭ�H��t�^a H��H�C(    �����H������H���   ����1ҋ�} ��b �e����H��t�a H�K8H�C0    ����H�Kh�;����:���fD  �����e���fD  H���X���H����������������S����UWVSH��H��(H�M(H�2} �����H�E(H�X8H��������=�O t����H�U(�} ��a ��` H�u(H�ىFp�R���H�E(H��H���   �'  ����   H��| ����H�E(H�X8H���{���H�E(H�H0H�pH��t�` H�E(H�x( H�@0    ��   H�������H���m���H�E(H�@8����ǀ�      H�a H�=Q| H����������   1�����H�4| ����H�E(H�@H����   H�}(H�O��H�Ð�H�| �����H�E(H���  H�XH���(����~�������H�E(H��� ﾭ��7���H������H�}( tH�E(H���   uH���b���1ҋ�{ ��` �8������;a ��   �t��� f.�     ��M �f�     UWVSH��8��M ��H�L$`H��tVH�D$`H��t\H�L$`����H�L$`H�h(�t����8��^ H�L$`���`���H�\$(A��A��H�l$ H�w� H���%  �H��8[^_]��    ��^ I��1�H�A� A��H��8[^_]�^%  @ f.�     1�� f.�     H��8�J^ H��H�T$ L�D$(�g^ �   ��t#H�T$ H��t1�H�Ѓ��H��u�ɸ   Dȉ�H��8�g       UWVSH��8�   H�-�] �ɉ�D�1���H�T$ H��L�D$(�^ ��t:H�D$ 1�H��t H�9�~�tH����H��u�H�D$     ��H��H����^ ��H��8[^_]�D  ATUWVSH��@�H��H��H��tk��t7����H�hH��H���p���D�#E��tZA��u"H�������H��tH������1�H��@[^_]A\ù   �y E��I��H��� H������뼸   H��@[^_]A\�H����H�|$(H�D$ �8���H��tCH�@H�D$0���"���H��tMH�T$ H�P�����
���H��t%H�T$0H�P�   �O����H�%    fD  H�D$0H�%    �H�D$ H�%    �AUATUWVSH��(�   H��H��H���#  H��x �d  �FK �DK 9�s=H��J ��L��I�8 ��   �QH�Љ��f�I��H��H�x� ��   ��9�u��t1L��J 1�I�8 I�@u��   I��H��H�x� ��   ��9�u��   ��   �ؽ   H�XJ D�c�AD�=   N�Hc�H������H��I����   ��A��1�M�L� A)�I��L���s���H��L�-	J H��w I����   HD�D�%EJ �-CJ I�9�  1�H��([^_]A\A]É�H���   �HD�H�Yw I�8�  1�H��([^_]A\A]�f�H�9w �d  �   �1��f�     WVSH�� �   9�I ����   H�=^I  ��   H��v ���  H�CI H�<�    9�I H��    v�}I H��v �y���H�JI H��t@H�FI H��H�H�H��t!L�BPM��t;ZHsI�8    H�H�RX�2 H��H9�u�H�^vh        �����H�Zv �  1�H�� [^_Ðf.�     UWVSH��(����Y ���)���H�xhH��H���z���9^Hv5H�FX�< t+H�FPH��H����������Z H��H��([^_]��    1���f�f.�     AWAVAUATUWVSH��(��I����Y A������H�hhH��H�������9sHv9H�{PL�4�H�CXH���0�!���D���Z 1�H��([^_]A\A]A^A_�D  H�KPD�fMc�J��    �����H��H��tSH�KXL�������H��I��t?�CHE��1�H��A)�I��������KHE��1�H��L�A)�����H�{PL�{XD�cH�X���H�������   �e����f.�     1�H9�����    H��u�f.�     �;����f.�     H��(����1�H��tH���  H��H��(ÐH��(�w���H��tH�@0H��(�f�     1���f�f.�     H��(����H��tH�@(H��(�f�     1���f�f.�     H��(����H�PH���    HE�H��(�f���F �1��D  1���F ��    VSH��8H�������H���  H�pH��ud�@@0uH���   �   �1  ��s �{X H��H��t1H�x( H�H0tqǀ�      H�ɋpt��V �CDH�C0    u���Y H�D$(�����H�D$(��ﾭ�H�K(��V H���   H�C(    t61ҋ+s �X �H��� ﾭ�t�~V H���   H�C0    �su�H���������f.�     H��(��E ��u1�H��(������H��H��t�@ ����B@t��BD�   t���@ SH�� ������H��tH�� ��~
�� H�� [���(H�� [� i       SH�� �f����   �P@H�Ã����P@������-E H�[H��tH�K�H�[H��u�1������ﾭ��;����f.�     SH�� �F���H��H��t�@@u���   ��u�CD����tH�� [�1�H�K0��V ��u�H�K8�$����O����@ f.�     VSH��(����H��H��t�@@u
�YD ��uH��([^�fD  H�s8H���4����C@�t<�SD��t4�K ��-H�K0��������SD�C@H��t��U H�����������f�H��H��([^����f�WVSH�� H��tt����H�ø����H9�v2����������H���@���H�O0H��tW����U �*���1�H�� [^_������H�ۉ�H��u�����1��pU �����1�H�� [^_�D  ������f�     ���DU �fD  VSH��(���s�����H��t,����H�N0H��t>���jU ����1�H��([^��     ����1���T �~���1�H��([^�D  ����T ��fD  UWVSH���  H���=���H��H����   H�H(H�A�H�����   H�l$ H����S ����   H�{8H���}�������1�H��tH���  H9��C@tE�SD����tf�u>������C@��IB H�K0H��t��S H�������1�H���  [^_]è��   H�������C@tܸ   H���  [^_]�D  �uبu�H�K(�D$P  ��S 1�H�K(�T =  u�H�K(H����R H����H�K(H��H��$  �~S �C@�cD�������C@���A H�K0H��t�>S H���
���H�K(��R �)���������C@��RA H�K0H��t�S �CDj       ������������H���CD�C@�����C@����������f�     VSH��(H�ˉ�H�&n �����H�������H��tMH9��  uD�@@u>���   ��u4H�@(H��H���w&H��m �I�����t5����w1H��H��([^����H��m �#����   H��([^��    1���   ��D  �!�Ðf.�     �   ��D��u	#1�D	�f.�     1�H�A    H�A    �A    �   H�A    H�A    �1�H�    H�A    H�A    H�A    �@ f.�     �   ������u����	�1����    ����1��fD  H��t�Ѓ��uD�A���D	��    �   �f.�     ����1��fD  �   ������u����	�1����    ����1��fD  H�AH�1��fD  1�H�Q�f�     H�AH�1��fD  1�H�Q�f�     UWVSH��(��H������H�ø   H��t������t	H��([^_]�H�k8H������H��t�CD����CDH���  ���	ƉsD�����H���(���1�H��([^_]� f.�     UWVSH��(��H������H�ø   H��t������t	H��([^_]�H�k8H���4���H��t�CD����CDH���  ���	ƉsD�@���H������1�H��([^_]� f.�     AVAUATUWVSH��@H��I��L��L������H��H���]  H��tH���  H�E L�%�O H�{H�=_N H�s1�ǃ�       �CD   H�C(����M��E1�E1�1ɺ   ��H��H�C0u)H��t�   A�փ�tH���А1�A����f�     k       H�shH�C8����H������H�{0 ��ǃ�       ǃ�       ��   1�M��tA�E A�U��CD�=  A�E���   1��D$    I��H�D$(    L�������O H��H�@�H���vcH�K0H��t�XM H�K8�����H������H�C0    H�C(    H��tH�E     H���   ��   �   H��@[^_]A\A]A^�@ ���   ��������| �����|���   ��   f.�     H���N H�K0��M �CDu'H�{(H����M 1���M 1�H��@[^_]A\A]A^ÐH��H�C(    �kM H���zL ��@ H�������K��� �T$<������T$<���   ���   ����f����   N��`���WVSH��@H��H�������H��H����   H�H(H����   H�T$<�NL ����   �CD�   ��   �n���1�H��tH���  H9���   ���   H�K(��t
H�A�H���w������HM H�K(H�5�K ��H�K0H��t��H��H�C0    tH�CH�H�K8�����H�Kh����1�H���   uH�ىD$,�����D$,��     �   H��@[^_� �$   ��f�     WVSH��0H��H��H��g �W���H���?���H��H����   H�H(H����   H�T$,�/K ����   �CD��   �T���1�H��tH���  H9���   ���   H�K(��u1��;L ��t���   ����   H�K(H�5~J ��H�K0H��t��H��H�C0    tH�CH�H�K8�����H�Kh����H���   t]H��f �!���1�H��0[^_��    H��f �����   H��0[^_��    H��f �l       �����   H��0[^_��    H�������fD  H�Qf �����$   �H�>f �����   �f.�     VSH��8�e���H�f H�������H����   H�K(H����   H�T$,��I ���}   �CD���   ��H�K(H�C(    �CDH��tBH�58I �֋��   ��t/H�K0H��t��H�K8H�C0    ����H�Kh�C���H���   tLH�ze �����1�H��8[^�@ H�ae ������   H��8[^��     H�Ae �����   ��H�������� ��7 �f�     1���7 ��    UWVSH��H�   H��H��H����   �/����   H��H����   H9��  ��   �@@��   ���   ����   H�@(H��H���w{H���C  H��H��t{H�N`H��t�����FpH�~`�D$    H�l$(�D$4    �D$0�{H ��u
H�=�6  tL�L$ A�   1ҹ�m@�}H ��H��H[^_]�fD  �   ��H��H[^_]û   ��f�     UWVSH��(�   H��H��H��L����   �,����   H����   H9��  ��   �@@��   ���   ����   H�P(H��H���w{H����   H�x`H����   H������H9�shH��H�����w[H��tf���u�]�H�Մ�tS�H�U�H��H��H��w�H��u:�F� �"   ��H��([^_]�fD  �   ��H��([^_]û"   ��f�     � �ʐ����������WVSH�� H��H�    H��H��b �@���H��tKH�H��tCH���t]�8�𱺾   u�p��u9H�H�    H��b �C�����H�� [^_�f�     m       �   ��f�     �   ��f�     H�    1��D  SH�� H��H�ib ����H��t:H��   H��t�8��uH����   t�@1�H�2b ������H�� [û   ��fD  WVSH�� H�yH��H����������t��H�� [^_�f.�     H�N ��������t�H��������H�� [^_�D  f.�     WVSH�� H�ˉ�H�I �����H�K���������t@��tH�� [^_�	�E�H�� [^_Ð1ҋA���A    �A� f.�     VSH��8H�ˉ�H�Fa ����H��8��u&H��@��~H�H�"a �h������H��8[^ù   ��` �D$ (   L�n� L��� H��H��� �����   �6���� f.�     �z3 �f�     UWVSH��X�b3 ��H��H��tKH�H��tP�h�8�1D H�H�t$@H��� A���D$0    H�D$8    �D$(    A���l$ ��
  �H��X[^_]�@ ��C H�I��H�o� A��H��X[^_]�
   f.�     ATUWVSH�� �   H��H��tzH�    �0   �   �   �N���H��H��tWH�h1�� ﰭ�H�@    H���@    �S�������uEL�f 1�L���?�������u)H�N(1���������u8���H�7��H�� [^_]A\�f�H���H���H��耼����H�� [^_]A\� H���(���L��� ���H���X����fD  SH�� H��H�!_ �l���H�;�tH�_ �   ������H�� [�1�H�������H��^ ���u�����H�� [� f.�     VSH��(H�9�H��tAH��^ �   � ���H�H��tn       �8��tH��^ �$�����H��([^Ã@1��� �K����������t���WVSH��0H��H�_^ ����H�T$(H���=���H�F^ ���������uHH�|$(H��t>H����������uC�G9G�G��~FH�D$(�   H��H��O����Å��   D؉�H��0[^_�f�     H�D$(H���H��0[^_�1��ﰭ�H����������u�H�O(�/���H�O����H�O �}���H�L$(�ﰭ�譺��또f.�     UWVSH��(H��������tH��([^_]� H�3H�~H��������u��F�~���tH��������H��H��([^_]�����D  H�N ���������tH���Y�������D  �F1��F    H��)F�9�����    UWVSH��(H��H���������t	H��([^_]�H�3H��H�nH��������u��F�~���tH���������H��H��([^_]�2���f�H�N H���T�������t=�   t'H���������ɋF1��F    H��)F�����f���F��f�     UWVSH��(H���P�����tH��([^_]� H�3H�~H��������u��F�~���tH���7�����H��H��([^_]����D  H�N �w�������tH���	�������D  �F1��F    H��)F�������    UWVSH��(H��������tH��([^_]� H�3H�~H���q�����uZH�N �d�������u>�F�   ��uA�V�F��~)��F    �F��~81�H���n����   ��D��H���X�����Dŉ�H��H��([^_]������F   1���D  WVSH��0H���a�����u]H�3�V��t#��n1�H��������H�o       �H��0[^_�S��� H�~ H���D�������u���F�F��t"H�����������fD  H��0[^_��     H�N(�w���H���D$,�����T$,��D��AUATUWVSH��HH���\�����tH��H[^_]A\A]�H�3H��� �������u&�V��u�V�F��~)��F    �F����F��H������H��H[^_]A\A]�H�t$(L�n �؉FH�H���H�D$ L�f(�z���H� H�D$0���j���H�T$ H�����F��y6L��L�����������t��@���H�T$0��H�H�L$(�T$ �t����     ����H�T$0H��F    �N����    AVAUATUWVSH��@H��H��H��t'H��t"�=�����t-H��@[^_]A\A]A^�f.�     �   H��@[^_]A\A]A^�H�;H��H�oH��������uVL�g H��L��������A��uP�W��u�W�G��~)��G    �G��O��GD��H���/����q���f.�     ��H�������X����H������D��H��������?����     H�|$(L�w(�؉GH�����H�D$ �����H� H�D$0�������H�T$ H����@ ��uEI��L��L�������ŋG��x�����H�T$0��H�tH�L$(A���T$ �9����G    �(�������H�T$0H����     H������fD  H��t1��    �f��   �f.�     H��tH��t��1�ø   �f�     H��t��w1��Ð�   Ð����������%6< ���%&< ���%< ���%< ���%�; ���%�; ���%�; ���%�; ���%�; ���%�; ���%�; ���%�; ���%f; ���%V; ���%F; ��p       �%6; ���%&; ���%; ���%; ���%�: ���%�: ���%�: ���%�: ���%�: ���%�: ���%�: ���%�: ���%v: ���%f: ���%V: ���%F: ���%6: ���%&: ���%: ���%: ���%�9 ���%�9 ���%�9 ���%�9 ���%�9 ���%�9 ���%�9 ���%~9 ���%n9 ���%^9 ���%N9 ���%>9 ���%.9 ���%9 ���%9 ���%�8 ���%�8 ��H�D$�H�G< � ��%v< ���%~; ���%f; ���%V; ���%�: ���%�: ��Ð��������������Ð��������������H��8I���I(�����tn��<tWv5L��    I��<u7I�RL�L$(MB��  H�D$(H��8�f.�     ��uL��    I����<t��>���fD  L�I����    E1�륐����������WVSH��0I� H�D$(H�H��H��L��H���P��tH�D$(H� H�D$(H�A�   H��H��L�D$(�P ��tH�T$(H�H��0[^_Ð��UWVSH��(1�H��H��H��L��t�#��H��H�w�����   H�C�H�V<��C(��   E1�1�D  H��D�B�L����H����I	�E��x�I�L�KH�B�E1�1ɈS)H��D�@�L��H���I	�E��x�I�L�K H��([^_]���H����   L�KI����H���R  H���H�V<��C(�c���H�C    뇐��UWVSH��(H�YI��H��H��L�D$`H�l$`L�1�1�f.�     H��D�C�L����H����H	�E��x�H��t#H�������I��H��H���H�����t�H��([^_]�1�H��([^_]�H��(���t/�ȃ�p< q       t>v<@t(<Pt<0u<H��H��(����@ ��t<u$1�H��(ÐH��H��(���@ H��H��(�����������������������SH�� ��w,��j�uH�B�H�Z@H��tH����H��H�� [�D H�� [�H�J��a  �VSH��(��PA��tR�����3  L�ߕ ��Ic�L��� M�I�@M��tD�ك�p��ID�I�E��x/M�H��([^�D  I�@H���L�H�@M�H��([^��    M�M�H��([^� L��E1�1��     H���p�H���H���I	�@��x��v���E�I�@�i���f�E�I�@�[���@ McI�@�K���@ L��E1�1��     H���p�H���H���I	�@��x��?������@�	���H������H��I	������M�I�@������F�����������������VSH��(���+���H���;@ ����H��H���KB H��H��t�M����@ ��������H��(���5 ������   ��= ������Ð��������������SH�� H��'	 H��H��� �   H��H�� [�= �������H��'	 H��q� ��   �f= ������Ð��������������SH�� H�$(	 H��H������   H��H�� [�'= �������H��'	 H������SH�� H�D(	 H��H��y����(   H��H�� [��< �������H�(	 H��Q����AWAVAUATUWVSH��   ��A��M��H�D$`    �D$\    ��   H� �Լ����I�0H��H�D$(�D$ �|$ ����@ ��D$C��   I�i�H���>  I�A�A�y�H�D$0��yPH�T$0L��$�   H��$   ������$�   Hr       ��$   �������$�   H��$   H��$�   �����I�E�H��$   M��1�� ��H��$   LcǺ   � ��H��$   H���D ���   ��   H�ĸ   [^_]A\A]A^A_�@ H��$   �# ��H��H�D$0�y  H�T$0H��$�   H��$   I��H�D$8�������$�   H��$   H������H��$   H�T$\H��$�   �����|$\H��H�� H;�$�   ��   L�d$hH�l$pH�|$x�     D��$�   1�D������I��M��D��H���\�����$�   1�I�ǉ�����M��I���H���8�����$�   1�I�ǉ��t�����I��M��H������E1�1�H��H���V�H�Ѓ�H����I	���x�H�D$hH�$�   H9�v_A��ty1�1�E1�H�|$(�   �����A�}�H�T$`H�|$0M�U�I�m�I�U�I�}��f���L����< H�l$xH��u?�   �J���f�HD$pH9�w�H9�$�   ������fD  A��uH�|$(v��- H�$�   M��u&H��t�A��u�D����uH�|$(�����1�����H��$�   H��N�T��x���M���  H��� H��D�����D$DuH�|$(H��� H����  �|$ H�l$ H�D$`I��D�d$CL��$  M�Ջl$DH�D$HD��$  L��E1�1� H���S�H�Ѓ�H����I	Ƅ�x��?w��@t�   H��H��I	�H��1�1�fD  D�H��L����H����H	�E��x��?wA��@t�   H��H��H	�M��tfl����@��t	M����   L��E1�1�H��H�$�   H��D�B�L����H����I	�E��x�M������uJH����   L�,3����D  s       A�   ��H�L$8L������H��tM��t�L�D$HL��H��������t�L��D��$  M��H�l$ L��$  A��������D$D��uH�|$(�u������������� �    L�D$`M��L��H�L$8��������H���E��H�l$ D��$  L��$  �i���D�����]���A��������_���f.�     A�E I�E@tI�E�H�D$`H��p���H�������H���U9 �N���SH�� ��L ��tH��v H�� [� H��L �$= ��t�H�iv 1��"���H�{L �V> H��A �*M��H�Cv H�� [�H�VL H���< H������������SH�� H�4"	 H��H��� H��H�� [�l6 ������������H�	"	 H��� ��K6 �����������Ð��������������H��(��K ��tH��u H��(�D  H��K �D< ��t�H��K �= H�MA �XL��H��u H��(Ð�������������5 �����������Ð��������������SH�� H��H�AN ��������%  H�5N L�K�H��tuL�[�O�L9�whH�J��   H����   I9�r�   f.�     I9�H��sH��H�AL�RH��u�I9�tSI�H�H�I9�t6H�@L�[�H�C�I�L�H�H�S�L��M H��M �������u[H�� [�I�L���fD  I�@MH�A� LH�K�L�[�L�fM �L�]M 1�H���s���L�LM H��H���a���H��#	 �   ��5 L�Q  H�H�W� H���= �  H��H��u�\7 ������������SH�� H��H��L 蜷������   H�K�   H�t       �L H��HB�H��H���H��t#L�L9�w�mD  L� L9�v(H��H�BH��u�1�H��L �޹����uNH��H�� [ÐH��M��L�PI)�I��vL�M�PH�M�H�L�H�X�f�L� L���H��H�6L ��H��"	 �   ��4 L�D  H�H�J� H���< �  H��H��u�O6 ����������������=��<��   H��� Hc�H���@ H��� ��     H�}� ��     H�q� ��     H�d� ��     H�[� ��     H�0� ��     H�7� ��     H�� ��     H��� ��     H��� ��     H�� ��     H�Ҋ ��     1�Ð������������H��Z H��Z ����H�'[ Ð�����H�)H H�H ����H�[ Ð�����ATUWVSH�� L�%K* ��H��L��L���
f�H)�t#H�A��H�������H�H���u�A�ԃ8t�H)�H��H�� [^_]A\Ð���������H��(H�	褷����uH��(ù   ��2 H�� 	 H�L�P  H��H�V� �: H��H��u�c4 �������������������H��H��� �������H��H�� ���������P �����������ATUWVSH�� H��H��D��H�sHM���j A��H��H��H��	 H��Y� H���1[  ��uH�� [^_]A\�f��{XH��L�cp�!O 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H����k H������������ATUWVSH�� H��M�̉�H�sHD����i A����H��H��	 H��� H���Z  ��uu       H�� [^_]A\�@ �{XH��L�cp�qN 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H���Mk H���5��������SH�� H���Si H�L	 H�H�� [Ð��ATUWVSH�� H��H��D��H�sHM���!i A��H��H��H�	 H���� H���Y  ��uH�� [^_]A\�f��{XH��L�cp�M 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H���}j H���e��������ATUWVSH�� H��M�̉�H�sHD���rh A����H��H�c	 H��� H���Y  ��uH�� [^_]A\�@ �{XH��L�cp��L 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H����i H�����������SH�� H����g H��	 H�H�� [Ð��SH�� H�D� H��H��H���O H�KH�<� H��� H�K8H��H��%� H��H�� [��- ��������SH�� H��� H��H��H��O H�KH��� H�U� H�K8H��H�H�� [��� SH�� H��� H��H��H��eO H�KH�� H�� H�K8H��H�H�� [�� H��H��� �������H��H�� ��������;p �����������ATUWVSH�� H��H��D��H�sHM���!� A��H��H��H�	 H��Y� H���1W  ��uH�� [^_]A\�f��{XH��L�cp�qn 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H��荋 H������������ATUWVSH�� H��M�̉�H�sHD���r� A����H��H�c	 H��� H��v       �V  ��uH�� [^_]A\�@ �{XH��L�cp��m 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H���݊ H���5��������SH�� H���ӈ H��	 H�H�� [Ð��ATUWVSH�� H��H��D��H�sHM��衈 A��H��H��H��	 H���� H���U  ��uH�� [^_]A\�f��{XH��L�cp��l 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H���� H���e��������ATUWVSH�� H��M�̉�H�sHD���� A����H��H��	 H��� H���U  ��uH�� [^_]A\�@ �{XH��L�cp�Al 1�H�C(    f�CyH�ChH�C     H�C0    H�CH�CH�CH�� [^_]A\�H��H���]� H�����������SH�� H���S� H�L	 H�H�� [Ð��SH�� H�T� H��H��H��Uo H�KH�<� H��� H�K8H��H��%� H��H�� [��) ��������SH�� H�� H��H��H��o H�KH��� H�e� H�K8H��H�H�� [��� SH�� H�Ļ H��H��H���n H�KH�� H�%� H�K8H��H�H�� [�� UATWVSH��H�� H��y I���������H�� H��L�d$ I�t$I���I��L��I��I��L��H��L��M�L)�I��	�A�w�L)�H9�wI)�I��I�T$�I�����H��[^_A\]ø���������ATUWVSH�� H��L��H��H�|��fD  �H��H�����ttH9���   <%u��V��st��ztt��%����H���fD  I�M�A���t)H��H)�H���    w       H9�toH��H���S����u�H���M����u�H��� H)�H�� [^_]A\��    �~u�V���M�M�aH��H��H)�������~H�H��M��H��6���H��H���  �H�A@Ð����������ATUWVSH��0H�AL�a8H��H�RH��H�|$(H�k8H�QH�SH�CH�AH�QH�SH�CH�AH�QH�S H�CH�A H�Q H�S(H�C H�A(H�Q(H�S0H�C(H�A0H�Q0L��H��H�C0�� H��L���� H��H���� H���J� H�F@H�S@H�V@�SHH�C@�FH�VH�CHH��0[^_]A\Ð��H�I@�ߖ���������SH�� H��H�I@�w����CHH�� [Ð�����VSH��(L�I@H��H�˺   H���k��������H��~�T��SHH��([^Ð���������L�I@H�к   H������������������VSH��8H��L��E1�H�����E��H���A    tE1�A��A��A��H�N@�����tH��H��8[^�D  H�N@����C    H�H��H��8[^Ð��VSH��HH��H��I�H�H�w���H�@ H9�uNH�N@E1�H������C    �����tH��H��H[^�fD  H�N@�G���C    H�H��H��H[^� D�L$ I��E1�H��H����H��H��H[^Ð��H��(��H�Q@���t��H��(鎔��fD  H���0�����������H��(Ð��������SH�� ���H�ˉ�u�KH���tH�S@������CH����H�� [� ���쐐����������SH�� H��H�I@�w���H�S@��H�� [�������������������VSH��(H��H���?R H�(	 H�H�C@H�F@�CH�FHH�C@    �CH����H��([^ÐVSH��(H�� H��H��H�Hx       ��H�A    H�I8H�A�    H�A�    H�A�    H�A�    H�A�    �� H��	 H�s@H��CH����H��([^ÐVSH��(H��H���Q H�x	 H�H�C@H�F@�CH�FHH�C@    �CH����H��([^ÐVSH��(H�S� H��H��H�H��H�A    H�I8H�A�    H�A�    H�A�    H�A�    H�A�    ��� H��	 H�s@H��CH����H��([^ÐSH�� H�� H��H�H��H�I8�a� H��H�� [�# ����H��� H��H�H��8�9� ���������VSH��(H��H���Q H�C@H�C@    H�F@�CH�CH�����FHH��H��([^Ð�������H�A@Ð����������ATUWVSH��0H�AL�a8H��H�RH��H�|$(H�k8H�QH�SH�CH�AH�QH�SH�CH�AH�QH�S H�CH�A H�Q H�S(H�C H�A(H�Q(H�S0H�C(H�A0H�Q0L��H��H�C0�� H��L���}� H��H���r� H���:� H�F@H�S@H�V@�SHH�C@�FHf�VHf�CHH��0[^_]A\Ð��������������H�I@鿑���������SH�� H��H�I@�G���f�CHH�� [Ð����UWVSH��(1�M��H��H��L��u�(fD  f�D] H��H9�t2H�N@����f���u�H��u1۸����f�FHH��H��([^_]��    �D]�f�FHH��H��([^_]Ð����������UWVSH��(1�M��H��H��L��u�#fD  H��H9�tH�W@�L] �)���f���u�H��H��([^_]Ð������VSH��8H��L��E1�H�����E��H���A    tE1�A��A��A��H�N@�������tH��H��8[^�D  H�N@�'���C    H�H��H��8[^Ð��y       VSH��HH��H��I�H�H�w���H�@ H9�uNH�N@E1�H������C    ������tH��H��H[^�fD  H�N@����C    H�H��H��H[^� D�L$ I��E1�H��H����H��H��H[^Ð��H��(H�A@f���t��H��H��(���� H��蠏����������H��(Ð��������SH�� f���H��u$�IH��f���t	H�S@�%��������f�SHH�� [����㐐�������SH�� H��H�I@�׎��H�S@��H�� [������������������VSH��(H��H���V H�	 H�H�C@H�F@�CHf�FH�����H�C@    f�CHH��([^Ð������������VSH��(H�s� H��H��H�H��H�A    H�I8H�A�    H�A�    H�A�    H�A�    H�A�    ��� H��	 H�s@H������f�CHH��([^Ð��������������VSH��(H��H����U H�H	 H�H�C@H�F@�CHf�FH�����H�C@    f�CHH��([^Ð������������VSH��(H��� H��H��H�H��H�A    H�I8H�A�    H�A�    H�A�    H�A�    H�A�    �� H��	 H�s@H������f�CHH��([^Ð��������������SH�� H�$� H��H�H��H�I8�� H��H�� [�D ����H��� H��H�H��8�i� ���������VSH��(H��H���U H�C@�����H�C@    H�F@�CHf�SHf�FHH��H��([^Ð���SH�� H�t	 H��H��y� H��H�� [� ������������H�I	 H��Q� �SH�� H�d	 H��H��9� �   H��H�� [� �������H�9	 H��� �SH�� H�z       T	 H��H���� H��H�� [�< ������������H�)	 H��Ѳ �UAWAVAUATWVSH��   H��$�   H�org/bugsI�gh spaceI� for forI�mat expaI�nsion (PH�lease suI�bmit fulI�l bug reI�port at I�https://H�/):
    H�M`H��H+u`H�not enouH�gcc.gnu.H�E�H�U�L�}�H�FxL�u�H���L�m�L�e�H�}�L�]�L�U�L�M�L�E�H�M�H�] �E ����H)�H�org/bugsH�T$ H�U`H�\$ L�D$hI��H�L$pH��$�   H�D$xH�/):
    L�|$(L�t$0L�l$8L�d$@H�|$HL�\$PL�T$XL�L$`H��$�   �/����D3h H���2� ��WVSH��0�=rZ  ��   �eZ � H����   H�XL�L$,1��;*�D$,������E1�1�H�H��������   H�5�, H���ֺ   A�0   H�r I�������T$,�   ��tC��H��H��������   ��A�   �   H�r I��踉���D$,��uH��踉����" ��H��H��趉��뻹   �	, A�-   �   H��q I���o����҉���   ��+ A�   �   H�Mq I���E���訉��H��H��ub� H�H���R�   H����I��A�   �   H��q �����   ��H��H�������   ��H�¹
   �����z �f����P �k �W���H���^ H���f���������SH�� H�	 H��H�良 �   H��H�� [�� �������H��	 H��a� �H��(�   � H�;	 H�L�����H��H�'� ��! ��H��(�   �� H��	 H�L�����H{       ��H�W� �! ��H��(H��0 H��t����H��0     H��(Ð����������H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����H�H9��Ð�����UWVSH��(H��H��L��D���g ��u#��wH�I��H��H��H�@(H��([^_]H�� H��([^_]Ð������VSH��(L��L��� ��tH�3H�C   �C   H��([^Ð�SH��@H�       H�D$(H�L��H�D$     L�L$ M� H�D$0    �P0�T$(1�����uH�D$ H��   H��@[Ð�������UWVSH��(H�\$pH;�$�   H��$�   H��D��t+L��H���p ��tH��o�G   1�H��([^_]�@ H�T$xL�L$h�A L�L$h��t�1��oH��([^_]Ð���������1�L9D$(���D�ÐUWVSH��(H��H��L��L���������u#H�MI��I��H��H�H�@0H��([^_]H��@ H��([^_]Ð������AWAVAUATUWVSH��(H��$�   L��$�   L��$�   H��$�   I��L��H��E��L���| ��uXL9���   H�NI��E��L��H�H��$�   L��$�   L��$�   H��$�   H�@8H��([^_]A\A]A^A_H���     M��H�] D�}x%L�1�I9����D��E1�H��([^_]A\A]A^A_�I���u��E   ��L��H���� ���]���D�}�Ő�����WVSH��0H�\$pL9�H��H��tH�NH��H�H�\$pH�@@H��0[^_H��L��L�D$(L�L$ �z L�L$ ��L�D$(tø   H��0[^_Ð��������������AWAVAUAT|       UWVSH��XL��I��H��$�   L���������A���?  D�oA����  H�D$0A�wM��H�D$ D����D$(�&@ H�H;D$0��  H���  �D$8	GH��H���e  I���D$8    I��D�l$<H�D$0    K�\>H�D$@    H��I�܃�A��u�T$(��t�E1�H��tI��I��H��tH�E N� I�K�L>L�L$ H��$�   H��P0��A���o���H�|$@u	����   �D$8��~M��u����D$8H�WH������H�D$0H�T$@H�H�D$8H�W��H�G~�tkA�F����D��H��X[^_]A\A]A^A_�H��H�L$@tH��tD�D$/� D�D$/��������G   �f.�     K�D>H�D$@�Q�����t�A�F������E�o�U���fD  �G��A���r���H�    �G   �_������������������AWAVAUATUWVSH��   H��$  L��$�   �CH��H��$�   D��$�   L��$�   t�A�CL;�$   �)  H��$�   H����  ����  H��$   �    �D$[ H+�$�   �D$ZH��$�    HI�E1�I��H�D$`H�D$H��$�   �u���D$T�   M����  I9��|  H��u��tl��D�k��  ��t
�C�z  E��E��uA�   A�   ��A���r  D�Ѓ�����  D��D������{��  A����  D�KA����  H��H���P  H��D�KH�D$`    H���D$p    D��$�   H�D$h    H�DD�L$tH��H���tM�$D�D$TI�L�M��tI9�A��D8T$Z��  �uH��$�   ��d  A���}       H�LH�|$HL��$�   H�H�T$ H�|$8H��$   H��$�   H�|$0H��$�   H�|$(�P8�|$p�ST$l�������A�щS��  E��L�H�L$`�n���M���n���H���������D�k�w���E��E��A���  ���F  D��1���~\��H�L$`��  ��A�����T$hH�E1��S�t���@ H��$�   H�H9�$   �?���A��A���}  A�    E!�A���  D�KA��H�    A�   �C   �4���D��H�Ĉ   [^_]A\A]A^A_�f.�     A�������������D$h	C�����@ �D$[�����fD  �T$hH��H�A�ƉS�����E��������E������D  ����   @����   ������������;���f.�     A��~A���@  �E�6  H��$�    H�L$`�����H��$�   ��  H��$�   D�T$\I��H��$   L��$�   H��$�   H� H��$�   H�|$ �P@D�T$\��A���3���f�     �E�I���H��$�    xKL�$�   L9�$   ��  ����  H��$�   H�H9�$   ��  A�   A�   �[��� H��$�   �D�\$\�o  H��$�   H��$   L��$�   H��$�   H� H�T$ H��$�   �P@D�\$\A��A���k���f�     D��������D  D��E��D����������$�   L�#H��$�    �C��   1�L�$�   L9�$   ��E1��D��C����H��$�   H���� ���������$�   E1��C�t���D  �t$Z�D$Z @ t$[�D$[��������N���H�T$`�{~       A��H��T$h�S�4���E1�H��$�   ��"����C   ����H�    A�   �C   �����E1��������A�   A�   �L��������������������������A�   �0����   A�   �   �1����������AVAUATUWVSH��0L��$�   M9�H��H��L��M����   D�vL��H��H��OD  H�F�t:H��H����H��tH���t%H�H�H�NL�M��H��H�L�d$ �P@��!I��H��M��u��   H��0[^_]A\A]A^�	�H��0[^_]A\A]A^�L����� �¸   ���`����ǐ��H�9i Ð�������WVSH��0H�qA��H���A H�1H�A    t-H�D$    L�i E1�1���� H��H��0[^_��     H�D$    L��h E1�1��� H��H��0[^_�H�H��H9�t�k
 H����������H��h Ð�������H��h Ð�������VSH��(H��D���?y��I������H��H�CH��H�tH���y��L�E1�H��H����� H��H��([^Ð����H�iK Ð�������H�)a Ð�������H�qK Ð�������H��` Ð��������   H�	H9�wH�A�H�AH9���Ð���WVSH�� H��H��H��L��� x��I��H��H��I��H�� [^_�    L�I�C�H��t?M��t:H��L9�IG�@ H��E�CtH��M��fD;tH��I��u�H��H���u��H������Ð������������H�L�J���������H������H�	L�I�M��tL�I9�IF� f;At
H��H���u�Ð��������������WVSH�� H��H��H��L���@w��I��H��H��I��H�� [^_�           SM��t5H�H�X�I9�s)H��F�@tH��M��fD;tH��I��u�I��I9�u�I������L��[Ð��������H�L�J������������  ��������H��Ð�����������H��(I��������H�L�H+P�L9�rH��(�L���f� ������WVSH�� H��H��H��L���`v��I��H��H��I��H�� [^_�    H������L�I�K�H��t/H�L9�IG�M��t H��E�CtH��M��fD;tH��I��u��H��H���u�Ð�H�L�J���������H������H�	L�I�M��tL�L9�IG���H��H���tf9At�Ð��������������WVSH�� H��H��H��L���u��I��H��H��I��H�� [^_�    SH�H�X�I9�sCJ�@M��tH��D�tH��M��fD9tH��I��u�L��[�fD  I��I9�tF�@��I�������ܐ������H�L�J���������H������H�	L�I�A��M9�s!fB;At
�!�fF9AuI��M9�u�H��������     L��Ð�����������H��(H�L�@�L9�s	H�PH��(�H�XL 諼 �����������H�H�P�H�PÐ����A��Ð���������A����Ð������H�H�P�H�DP�Ð��H�H�P�H�PÐ���SH�� I��H�L��H�Z�I9�w>L)�L9�IG�H��tJ�JH��tL�L����t��H��H�� [��fA�H��H�� [�H��K I��I��H�WK �� ��H�Ð�����������WVSH�� H��H��H��L���s��I��H��H��I��H�� [^_�    WVSH�1M��L�^���   M9�H������vHN�FL��L)�I9�w9�   L)�M��H�t!H��t�
J�<^M�Y��fA;
tI��       �H��u�H������[^_�D  L9�tM1�L9�tFE�DBH��fD;Bt�I��H��L)�H��I9�w�H�M��t�H��u��f�M9�H������IC�[^_�L��H)�H��뚐��H�L�J��$�������H������L�	I�I�I9�s$L)�O�AM��t�fA9tI��H��u�H��������     M)�L��H��Ð�����H�H��H�Ð�����H�H�@�Ð�������H�Ð�����������H�Ð�����������H�H��H�Ð�����H�H�x� ��Ð���H�Ð�����������WVSH�� H��H��H��L����q��I��H��H��I��H�� [^_�    H������L�I�J�I9�wTM�Y�L)�L��L9�HF�M�BM��t:I9�t5M��A��H����A8�u,�
fA9u#1��E�THH��fD;JuI9�u���     H�H�I��H��tH���H������Ð�����H�L�J��d�������H������H�	L�I�M��tL�L9�IG� f9At
H��H���u�Ð��������������H�H��Ð�������H�Ð�����������H�H�@�Ð�������H�H��H�J�H�JH�Ð�������������SH�� H�H�@�H��I9�w�' H��H�� [�H��I I��H��G �h� ��������H�Ð�����������H�H�P�H�PÐ���WVSH�� H�H�X�H��H��H���p��H9�H��HF�H��tUL�L9�tMM��A��H����A8�tH�������H�� [^_��    1��<NfA9<HuCH��H9�u�f.�     H)ø���H������@H��   �M�H�� [^_�f.�     ���H�� [^_Ð��L�	L�I�A�I�H�I��H9�LF�M��t#M9�t1�E�PfE9Qu2�       H��L9�u��    H)�H�¸���H������@H��   �M�����Ð�������UWVSH��(H�H�X�H��H��L��H9���   H)�L��L9�IG���n��H9�H��HF�H��t^H�U L�zI9�tQM��A��H����A8�tH�������H��([^_]�f.�     1��<VfA9<PuCH��H9�u�f.�     H)ø���H������@H��   �M�H��([^_]�f�     ���H��([^_]�H��E I��I��H�F �� ���������H��(L�L�T$PI�C�H9���   H)�L��L9�LF�M9�IF�H��tNI�SL9�tEH��A��M����A8�tI�������H��(�f�1�E�AfD9Bu6H��H9�u�f�     M)и���I������@I��   �AM�H��(����H��(�H��D I��I��H�ME �I� ���������H��(L�I�C�H9�w~M�	H)�L9�LF�I�I�M��L9�LF�M��t0I�SL9�t'H�Ҹ����t<1�E�AfD9Bu3H��L9�u�fD  I)ȸ���I������@I��   �AM�H��(����H��(�H�D I��I��H��D 虴 ���������VSH��(H�L�T$`L�\$hH�C�H9���   I�1L�N�M9���   H)�L9�LF�M)�M9�MG�L��M9�IF�H��tQN�VH�SI9�tDH��A��M����A8�tI�������H��([^�1�f�     A�4Bf94Bu5H��H9�u�M)ȸ���I������@I��   �AM�H��([^�fD  ���H��([^�H�C I��I��H��C 蛳 H��C M��H��B 腳 �����H�H��H�J�H�JH�Ð�������������H��(H�	L�       �I�H��L��I9�rH��(�H��B I���6� ������H�H�@�H)�L9�IG�Ð�������������H�H�@�Ð�������H��������Ð����H�Ð�����������H�H�PÐ�������H�AÐ�����������Ð������������Ð������������   H�	H9�w
HI�H9���Ð�������WVSH�� H��H��H��L���j��I��H��H��I��H�� [^_�    UWVSH��(H�1H�F�H��L��H��tFM��tAH��L��L9�HF���H��H���t�I��H����j��H��t�H��H��([^_]�fD  H������H��H��([^_]Ð������������H�L�J��t�������H������H�	L�I�M��tL�I9�IF� :t
H��H���u��WVSH�� H��H��H��L���i��I��H��H��I��H�� [^_�    ATUWVSH�� M��I��L��L��tHH�9H�o�I9�r�:f.�     H��H9�t'�I��L����i��H��t�H��H�� [^_]A\�D  H������H�� [^_]A\Ð�������������H�L�J��t����������8  ��������H��Ð�����������H��(I��������?H�L�H+P�L9�rH��(�L���V� ������WVSH�� H��H��H��L���h��I��H��H��I��H�� [^_�    UWVSH��(H������H�9H�G�H��L��H��t-H�L9�IG�H��t�I��H����h��H��t
H��H���u�H��H��([^_]Ð�����H�L�J���������H������H�	L�I�M��tL�L9�IG���H��H���t8t��WVSH�� H��H��H��L����g��I��H��H��I��H�� [^_�    ATUWVSH�� H�1H�n�I��L��L��I9�sAM�       ��u�'f.�     H��H9�t'�I��L����g��H��u�H��H�� [^_]A\�D  H������H�� [^_]A\Ð�������������H�L�J��t�������H������H�	L�I�A��M9�s B:t
�"f�F8uI��M9�u�H�������f�     L��Ð�����������H��(H�L�@�L9�sH�H��(�H�	< �|� ������������H�H@�Ð��������A��Ð���������A����Ð������H�H�P�H�D�Ð��H�H@�Ð�������SH�� H�H�X�I��L��I9�w;L)�L9�IG�H��tH�H��tI��L���f��H��H�� [��A�H��H�� [�H�; I��I��H��; 赭 �����H�Ð�����������WVSH�� H��H��H��L����e��I��H��H��I��H�� [^_�    AVAUATUWVSH�� H�9M��H��L��H�W��}   L9�H������vbH�,L)�J�I9�wRA�   M)�L�I��tAD�.D����e��H��I��t&I��H��H���e����tII�NI��I)�L9�wM�u�H������H�� [^_]A\A]A^�L9�H������IC�H�� [^_]A\A]A^�f�L��H)��ʐ�������H�L�J��$�������VSH��(H������H�1H�F�I9�sJ�L)���I���%e��H��H)�H��HE�H��H��([^Ð�������������H�H��H�Ð�����H�H�@�Ð�������H�Ð�����������H�Ð�����������H�H��H�Ð�����H�H�x� ��Ð���H�Ð�����������WVSH�� H��H��H��L����c��I��H��H��I��H�� [^_�    UWVSH��(H������H�9H�G�H��L��I9�w6L)�L��L9�HF�H��t$H�I�       ��H���d����tH�C�H��tH��H��u�H��H��([^_]�H�������됐��H�L�J���������H������H�	L�I�M��tL�L9�IG� 8t
H��H���u��H�H��Ð�������H�Ð�����������H�H�@�Ð�������H�HR�H��H�Ð�SH�� H�H�@�H��I9�w��� H��H�� [�H�t9 I��H��7 �x� ��������H�Ð�����������H�H@�Ð�������UWVSH��(H�9H�_�H��H���vb��H��H9�I��LF�M��tH��H����b����uH)����H������@H��   �M�H��([^_]Ð�������������VSH��(H�	H�H�Y�H�r�I��H9�LF�M��t	�pb����uH)����H������@H��   �M�H��([^Ð��������������ATUWVSH�� H�1H�^�H��M��H9�w]H)�L��L9�IG��a��H9�I��H��LF�M��tH�.L����a����uH)�����H������@H��   �M�H�� [^_]A\�H�P6 I��I��H��6 �� ��������������VSH��(H�	H�t$`H�Y�H9�wMH)�L9�IG�I��H9�LF�M��tH�L���]a����uH)����H������@H��   �M�H��([^�H��5 I��I��H�G6 �c� ���VSH��(H�	H�Y�H��H9�wQH)�I�L9�IG�H�r�I��H9�LF�M��tH���`����uH)����H������@H��   �M�H��([^�H�C5 I��I��H��5 �� �VSH��(H�	L�T$`L�\$hH�Y�H9�wfI�H�p�I9�wsH)�L9�IG�L)�L9�IG�I��H9�LF�M��tL�H�H���?`����uH)����H������@�       H��   �M�H��([^�H��4 I��I��H�)5 �E� H�5 I��M��H��4 �,� ������������H�HR�H��H�Ð�H��(H�	L�I�H��L��I9�rH��(�H�>4 I���� ������H�H�@�H)�L9�IG�Ð�������������H�H�@�Ð�������H��������?Ð����H�Ð�����������H�H�Ð��������H��E Ð�������H��(H��H�JL�M�H(D�H��R  I9�uD� H�HH��(� H��H�D$0H��A��H�D$0H��(Ð�������H�9  H�H�@PH9�uH�A�@`�D  H���������������H�  H�H�@HH9�uH�A�@\�D  H���������������SH��0H�H�@(H��H��  H9�u%H�BL�D$/H��H�P(�z H��H��0[��    H����H��H��0[Ð�SH��0H�BH�PL�D$/H���vz H��H��0[Ð������������H�y  H�H�@@H9�uH�A�@X�D  H���������������H�Y  H�H�@H9�uH�A�@!�@ H���������������H�A�@`Ð�������H�A�@\Ð�������SH��0H�H�@8H��H�
  H9�u%H�BL�D$/H��H�PH�y H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H��   H9�u%H�BL�D$/H��H�P8�`y H��H��0[��    H����H��H��0[Ð�H��   H�H�@H9�uH�A�@"�@ H���������������SH��0H�BH�P(L�D$/H����x H��H��0[Ð������������H�A�@XÐ�������H�A�@!Ð������SH��0H�BH�PHL�D$/H���x H��H��0[Ð�����       ��������SH��0H�BH�P8L�D$/H���vx H��H��0[Ð������������H�A�@"Ð������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P� x H��H��0[��    H����H��H��0[Ð�H�9  H�H�@PH9�uH�A�@`�D  H���������������H�  H�H�@HH9�uH�A�@\�D  H���������������SH��0H�H�@(H��H��  H9�u%H�BL�D$/H��H�P(�pw H��H��0[��    H����H��H��0[Ð�SH��0H�BH�PL�D$/H���6w H��H��0[Ð������������H�y  H�H�@@H9�uH�A�@X�D  H���������������H�Y  H�H�@H9�uH�A�@!�@ H���������������H�A�@`Ð�������H�A�@\Ð�������SH��0H�H�@8H��H�
  H9�u%H�BL�D$/H��H�PH�pv H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H��   H9�u%H�BL�D$/H��H�P8� v H��H��0[��    H����H��H��0[Ð�H��   H�H�@H9�uH�A�@"�@ H���������������SH��0H�BH�P(L�D$/H���u H��H��0[Ð������������H�A�@XÐ�������H�A�@!Ð������SH��0H�BH�PHL�D$/H���fu H��H��0[Ð������������SH��0H�BH�P8L�D$/H���6u H��H��0[Ð������������H�A�@"Ð������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P��t H��H��0[��    H����H��H��0[Ð�H�9  H�H�@PH9�uH�A�@`�D  �       H���������������H�  H�H�@HH9�uH�A�@\�D  H���������������SH��0H�H�@(H��H��  H9�u%H�BL�D$/H��H�P(�P� H��H��0[��    H����H��H��0[Ð�SH��0H�BH�PL�D$/H����s H��H��0[Ð������������H�y  H�H�@@H9�uH�A�@X�D  H���������������H�Y  H�H�@H9�uH�A�@"�@ H���������������H�A�@`Ð�������H�A�@\Ð�������SH��0H�H�@8H��H�
  H9�u%H�BL�D$/H��H�PH�P� H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H��   H9�u%H�BL�D$/H��H�P8� � H��H��0[��    H����H��H��0[Ð�H��   H�H�@H9�uH�A�@$�@ H���������������SH��0H�BH�P(L�D$/H���� H��H��0[Ð������������H�A�@XÐ�������H�A�@"Ð������SH��0H�BH�PHL�D$/H���F� H��H��0[Ð������������SH��0H�BH�P8L�D$/H���� H��H��0[Ð������������H�A�@$Ð������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P�q H��H��0[��    H����H��H��0[Ð�H�9  H�H�@PH9�uH�A�@`�D  H���������������H�  H�H�@HH9�uH�A�@\�D  H���������������SH��0H�H�@(H��H��  H9�u%H�BL�D$/H��H�P(�� H��H��0[��    H����H��H��0[Ð�SH��0H�BH�PL�D$/H���p H��H��0[Ð�����       ��������H�y  H�H�@@H9�uH�A�@X�D  H���������������H�Y  H�H�@H9�uH�A�@"�@ H���������������H�A�@`Ð�������H�A�@\Ð�������SH��0H�H�@8H��H�
  H9�u%H�BL�D$/H��H�PH�� H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H��   H9�u%H�BL�D$/H��H�P8��� H��H��0[��    H����H��H��0[Ð�H��   H�H�@H9�uH�A�@$�@ H���������������SH��0H�BH�P(L�D$/H���V� H��H��0[Ð������������H�A�@XÐ�������H�A�@"Ð������SH��0H�BH�PHL�D$/H���� H��H��0[Ð������������SH��0H�BH�P8L�D$/H����� H��H��0[Ð������������H�A�@$Ð������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P�`n H��H��0[��    H����H��H��0[Ð�Ð��������������H�AH�HH�
H�@H�BÐ�����������H�AH�H H�
H�@(H�BÐ�����������H�AH���   H�
H���   H�JH���   H�JH���   H�JH���   H�J H���   H�J(H���   H�B0Ð��������������H�AH�H0H�
H�@8H�BÐ�����������H�AH��(  H�
H��0  H�JH��8  H�JH��@  H�JH��H  H�J H��P  H�J(H��X  H�J0H��`  H�J8H��h  H�J@H��p  H�JHH��x  H�JPH���  H�BXÐ�������AVAUATUWVSH�� I��H��1�1�M��M���P��H��H����O��H��       XH����� I��H��H��H���%P��I�V 1���O��M��L��H��L��$�   �O��1�H��H����O��H���o� H��u�E  H�� [^_]A\A]A^�H��H��t�ɧ���T� ����H�AH�HXH�
H�H`H�JH�HhH�JH�HpH�JH�HxH�J H���   H�J(H���   H�B0Ð�������������H�AH�H@H�
H�@HH�BÐ�����������H�AH���   H�
H���   H�JH���   H�JH���   H�JH���   H�J H���   H�J(H���   H�J0H��   H�J8H��  H�J@H��  H�JHH��  H�JPH��   H�BXÐ�������Ð��������������H�AH�HH�
H�@H�BÐ�����������H�AH�H H�
H�@(H�BÐ�����������H�AH���   H�
H���   H�JH���   H�JH���   H�JH���   H�J H���   H�J(H���   H�B0Ð��������������H�AH�H0H�
H�@8H�BÐ�����������H�AH��(  H�
H��0  H�JH��8  H�JH��@  H�JH��H  H�J H��P  H�J(H��X  H�J0H��`  H�J8H��h  H�J@H��p  H�JHH��x  H�JPH���  H�BXÐ�������AVAUATUWVSH�� I��H��1�1�M��M���M��H��H����L��H�XH����� I��H��H��H���M��I�V 1���L��M��L��H��L��$�   �4L��1�H��H���L��H���_� H��u1�f�E H�� [^_]A\A]A^�H��H��t跤���B� ��H�AH�HXH�
H�H`H�JH�HhH�JH�HpH�JH�HxH�J H���   H�J(H���   H�B0Ð�������������H�AH�H@H�
H�@HH�BÐ����       ��������H�AH���   H�
H���   H�JH���   H�JH���   H�JH���   H�J H���   H�J(H���   H�J0H��   H�J8H��  H�J@H��  H�JHH��  H�JPH��   H�BXÐ�������UWVSH��(H�� H����G  H��H�H�@H�<�H�H��tH��([^_]�f.�     ��   �6� H���@    H��H��n H�C    H��H�C    �C  H��H�C(    H�1�H�C0    H�C8    H�C@    f�CHƃ�    ��$ H�I��H���{ H�H��([^_]�H���� �[� H���� H�H���P��H���� H��踢����������UWVSH��(H�� H����F  H��H�H�@H�<�H�H��tH��([^_]�f.�     ��   �6� H���@    H��H��m H�C    H��H�C    �C  H��H�C(    H�H�C0    H�C8    H�C@    �CH    ƃ�    �q) H�I��H���z H�H��([^_]�H���� �Z� H���� H�H���P��H���� H��跡���������UWVSH��(H��
 H����E  H��H�H�@H�<�H�H��tH��([^_]�f.�     �p   �6� H���@    H��H�"� H�C    H��H�1�H�C    f�C �C" H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co �F H�I��H���ly H�H��([^_]�H���� �C� H���� H�H���P��H���� H��蠠������������������UWVSH��(H��	 H���D  H��H�H�@H�<�H�H��tH��([^_]�f.�     �       �p   �� H���@    H��H�"� H�C    H��H�1�H�C    f�C �C" H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co �JL H�I��H���Lx H�H��([^_]�H���x� �#� H���k� H�H���P��H���x� H��耟������������������UWVSH��(H�� H���C  H��H�H�@H�<�H�H��tH��([^_]�f.�     ��   ��� H���@    H��H�"� H�C    H��H�H�C    �C  �C"    H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz ��Q H�I��H���+w H�H��([^_]�H���W� �� H���J� H�H���P��H���W� H���_������������������UWVSH��(H�q H���iB  H��H�H�@H�<�H�H��tH��([^_]�f.�     ��   ��� H���@    H��H�"� H�C    H��H�H�C    �C  �C"    H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz �)X H�I��H���v H�H��([^_]�H���7� ��� H���*� H�H���P��H���7� H���?������������������H�AÐ����������H�9 ��Ð�������H��8H�AH�L$`L�L$ M��I��H��H�L$(1��� H��8Ð���H��8H�AH�L$`L�L$ M��I��H��H�L$(1��Y� H��8Ð���VSH��xH�RH�t$@H��1�L�L$ H�D$`    M��I���C� H�|$` t0L�D$HL�L$?H��H�T$@�$a H�D$`H��tH��       ���H��H��x[^�H�� �O� H�T$`H��H��tH����H���%��������VSH��hH�RH�t$0H��1�L�L$ H�D$P    M��I���� H�|$P t8H�T$0H�CE1�H��L�D$8H�I��\� H�D$PH��tH����H��H��h[^�H�l 跃 H�T$PH��H��tH����H��荛���������������H��8H�AH�L$`L�L$ M��I��H��H�L$(1��Y� H��8Ð���H��8H�AH�L$`L�L$ M��I��H��H�L$(1��	� H��8Ð���VSH��xH�RH�t$@H��1�L�L$ H�D$`    M��I����� H�|$` t0L�D$HL�L$?H��H�T$@�� H�D$`H��tH����H��H��x[^�H�T 迂 H�T$`H��H��tH����H��蕚�������VSH��hH�RH�t$0H��1�L�L$ H�D$P    M��I����� H�|$P t9H�CH�T$0E1�H��H�H�D$8L�B�� H�D$PH��tH����H��H��h[^�H�� �&� H�T$PH��H��tH����H�������������������VSH��xH��$�   H�R H�t$@H��H�HH�D$`    H�L$8H� 1�D�L$ E��I��H�D$0��$�   �D$(�� H�|$` t8H�T$@H�CE1�H��L�D$HH�I��� H�D$`H��tH����H��H��x[^�H� �c� H�T$`H��H��tH����H���9������������VSH��   H��$�   H�R H� H��H�D$p    H�t$PH�H�H�D$0��$�   D�L$ E��I��H�L$81ɉD$(��� H�|$p t3L�D$XL�L$OH��H�T$P�}] H�D$pH��tH����H��H�Ĉ   [^�H�: 襀 H�T$pH��H��tH����H���{��������������H��8H��H�Q L�D$ �       1�L�HL� �� H��8Ð������������H��8H�H�Q 1�L�H�L�D$ I����� H��8Ð������������A��H�Q 1��r� ��A��H�Q 1��R� ��VSH��xH��$�   H�R H�t$@H��H�HH�D$`    H�L$8H� 1�D�L$ E��I��H�D$0��$�   �D$(�� H�|$` t9H�CH�T$@E1�H��H�H�D$HL�B�W� H�D$`H��tH����H��H��x[^�H� �b H�T$`H��H��tH����H���8�����������VSH��   H��$�   H�R H� H��H�D$p    H�t$PH�H�H�D$0��$�   D�L$ E��I��H�L$81ɉD$(�� H�|$p t3L�D$XL�L$OH��H�T$P�� H�D$pH��tH����H��H�Ĉ   [^�H�: �~ H�T$pH��H��tH����H���{��������������H��8H��H�Q L�D$ 1�L�HL� �� H��8Ð������������H��8H�H�Q 1�L�H�L�D$ I���� H��8Ð������������A��H�Q 1��� ��A��H�Q 1��r� ��SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@d   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�軝 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@d   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�軛 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@t   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��ۜ H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@t   L�L$`)D$�       P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��ۚ H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@y   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1���� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@y   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1���� H��H��p[Ð�H�Q1���� �����H�Q1���� �����SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@w   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1���� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@w   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1���� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@m   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@m   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@d   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��[� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@d   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��[� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�       �   H���D$@t   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��{� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@t   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1��{� H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@y   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�蛚 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@y   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�蛘 H��H��p[Ð�H�Q1��� �����H�Q1��u� �����SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@w   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�蛙 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@w   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�蛗 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@m   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�軘 H��H��p[Ð�SH��pH��$�   �Ao�AoH�D$8H��$�   H���D$@m   L�L$`)D$P)L$`H�D$0H��$�   H�D$(H�D$PH�D$ L�B1�軖 H��H��p[Ð�AUATUWVSH���   I�0I�X�AoH��$X  H��$�   H��)D$PH�D$8H��$H  H�L$pL��$�   H�D$@    L�d$HL�L$`HǄ$�       H�D$0��$@ �        Ǆ$�       H�t$`H�\$h�D$(H�D$PH�D$ L�B1��)� H�    �����D$xH!Ӌ�$�   H�t$pH	�H��$�   ��t.H��$P  �H��H�7H�_tL����H��H���   [^_]A\A]�H����   H��$�   L��$�   E1�L��$�   I�EL��H��$�   I��D� H��$�   I�MH�E L�EH9���   L9�L��$�   H��$�   tWH��L�EH�U L�MH�MtNH��$�   L��$�   HǄ$�       I���  H��$�   L9�t��� H��$�   ����H�U L�MH�MI�EH��$�   봐L��H���5� H��$�   �H�� ��r H��$�   H��H��tL����H���Ҋ����AUATUWVSH���   I�0I�X�AoH��$�   H��)D$PH�D$8H��$(  H�L$pH��$�   H�D$@    H�l$HL�L$`HǄ$�       H�D$0��$   Ǆ$�       H�t$`H�\$h�D$(H�D$PH�D$ L�B1��� H�    �����D$xH!Ӌ�$�   H�t$pH	�H��$�   ��t5H��$0  �H��H�7H�_tH����H��H���   [^_]A\A]��    H��tlL��$�   L��$�   H��$�   L��$�   M��L���`N H��$8  L���`< H��$�   �������A���~H��$�   �r���H��L���!: ��H�� �cq H���H��H��$�   L��H�H��: H��$�   H��tH����H�������������������VSH��   I� I�X�AoH�D$`H��$�   H��H�D$@H��$�   H�D$8H��$�   H�L$pH�D$H    L�L$`H�\$h)D$PH�D$0��$�   Ǆ$�       �D$(H�D$PH�D$ L�B1��3� �T$�       xH�    ����H!�H�D$pH	Ӌ�$�   ��u/H��$�   ۬$�   �:H�H��H�^H�Ĩ   [^�f.�     H��$�   ��֐���VSH��   I� I�X�AoH�D$`H��$�   H��H�D$@H��$�   H�D$8H��$�   H�L$pH�D$H    L�L$`H�\$h)D$PH�D$0��$�   Ǆ$�       �D$(H�D$PH�D$ L�B1��s� �T$xH�    ����H!�H�D$pH	Ӌ�$�   ��u/H��$�   ۬$�   �:H�H��H�^H�Ĩ   [^�f.�     H��$�   ��֐���UWVSH��  )�$�   �Ao �Ao	H��$h  H��$�   H��)D$PH�D$8H��$X  H��$�   H�|$HH��$�   H�D$@    L�L$p)L$`H�D$0��$P  HǄ$�       Ǆ$�       )D$p�D$(H�D$`H�D$ L�B1��� ��$�   H��$�   ��H�D$PH��$�   fot$PfĴ$�   t4H��$`  �H��3tH���А(�$�   H��H��  [^_]�D  H����   H��$�   H��$�   E1�H�EH��H��$�   H��$�   L�B�ķ H��$�   H�UH�L�FH9�t|L9�H��$�   L��$�   tWH��L�FH�L�NH�Vt/H��$�   L��$�   H��1�HǄ$�       H9�f�t�� H��$�   �����    H�L�NH�V�� H��H����� H��$�   �H�� �?m H��$�   H��H��tH����H��������UWVSH���   )�$�   �Ao �Ao	H��$�   H��)D$PH�D$8H��$8  H��$�   H�t$HH��$�   H�D$@    L�L$p)L$`H�D$0��$0  HǄ$�       Ǆ$�       )�       D$p�D$(H�D$`H�D$ L�B1�輖 ��$�   H��$�   ��H�D$PH��$�   fot$PfĴ$�   t/H��$@  �H��3tH���А(�$�   H��H���   [^_]�H��tvL��$�   H��$�   H��$�   H��$�   I��H���� H��$H  H���Ͳ H��$�   �������A���~H��$�   �x���f.�     H��H���D� ��H�+� �k H���H��H��$�   H��H�H��*� H��$�   H��tH����H���P�������������������SH��   �Ao�AoH��$�   H��)L$PH�D$@H��$�   H�D$8H��$�   L�L$pH��$�   )T$`H�D$H    Ǆ$�       H�D$0��$�   )L$p�D$(H�D$`H�D$ L�B1��� H��$�   H�D$P��$�   foD$PfĄ$�   ��u H��$�   ۬$�   �8H��H�İ   [�H��$�   �H��H�İ   [Ð�SH��   �Ao�AoH��$�   H��)L$PH�D$@H��$�   H�D$8H��$�   L�L$pH��$�   )T$`H�D$H    Ǆ$�       H�D$0��$�   )L$p�D$(H�D$`H�D$ L�B1��#� H��$�   H�D$P��$�   foD$PfĄ$�   ��u H��$�   ۬$�   �8H��H�İ   [�H��$�   �H��H�İ   [Ð�ATUWVSH��   )�$�   H��$  �Ao8D��$  H�\$pH��L�@H��H�SD��H��HǄ$�       H�T$pH�E1�I��N� H�W� L�E1�H����E��@��H�\$@H��$�   H�D$PH�D$8H��$   L�L$`D�d$0�t$ )|$`H�D$(�|$P�Ĕ H��$�   H��tH���А�       (�$�   H��H�İ   [^_]A\�H��$�   H��H��tH����H���[��������������AUATUWVSH��   )�$�   H��$   �Ao8��$  H�\$pI��I��HǄ$�       H��H��D���E H�@��@��1�M�E��L��L�L$`H�@�H�\$@�l$0�|$ )|$`H�D$xH�� H��$�   H�D$PH�D$8H��$  �|$PH�D$(�� H��$�   H��tH���А(�$�   L��H�ĸ   [^_]A\A]�H��$�   H��H��tH����H���P������������������SH��pH��$�   �Ao �(E��H��)D$`D�L$ H�D$@    H�D$PH�D$8��$�   L�L$`�|$P�D$0H��$�   H�D$(L�B1��K� H��H��p[Ð�SH��pH��$�   �Ao �(E��H��)D$`D�L$ H�D$@    H�D$PH�D$8��$�   L�L$`�|$P�D$0H��$�   H�D$(L�B1�苒 H��H��p[Ð�ATUWVSH��   )�$�   H��$  �Ao8��$  H�\$pI��H��HǄ$�       H�SD��H��H�T$pH�E1�H�@L�B莰 M�D$��@��1�H��� H�\$@H��H��$�   H�D$PH�D$8H��$   ��|$0L�L$`�t$ )|$`H�D$(�|$P�e� H��$�   H��tH���А(�$�   H��H�İ   [^_]A\�H��$�   H��H��tH����H���\}��������������AUATUWVSH��   )�$�   H��$   �Ao8��$  H�\$pI��I��HǄ$�       H��H��D���P� H���@��1�M�E��L��L�L$`H�@�H�\$@�l$0�|$ )|$`H�D$xH�D� H��$�   H�D$PH�D$8H��$  �|$PH�D$(謔 H��$�       �   H��tH���А(�$�   L��H�ĸ   [^_]A\A]�H��$�   H��H��tH����H���Q|���SH��pH��$�   �Ao �(E��H��)D$`D�L$ H�D$@    H�D$PH�D$8��$�   L�L$`�|$P�D$0H��$�   H�D$(L�B1���� H��H��p[Ð�SH��pH��$�   �Ao �(E��H��)D$`D�L$ H�D$@    H�D$PH�D$8��$�   L�L$`�|$P�D$0H��$�   H�D$(L�B1��;� H��H��p[Ð�H�h
 Ð�������H��H�7����������H��H�'����������H�AÐ����������H��`�����������H�AÐ����������H��`������������H�AÐ�����������Ð������������Ð�����������H�AÐ����������H�AÐ����������H��X�����������H�AÐ����������H��X�g����������H�AÐ����������H��P�G����������H�AÐ����������H��P�'����������H�AÐ����������H�A(Ð����������H�AÐ����������H�AÐ����������H�A0Ð����������H�A Ð����������SH�� H��H��8��m H��H�� [Ð�����H�AÐ����������H�A(Ð����������H�AÐ����������H�AÐ����������H�A0Ð����������H�A Ð����������SH�� H��H��8�Om H��H�� [Ð������A����������Ð�������������H��HH�T$xH��H�T$0H��$�   L�D$ D�@H�L$ L�L$(D�HH�T$8H�T$0��n H�T$pH�L$ H�
H��$�   H�L$0H�
H��HÐ��������������VSH��8H�D$x�A��       YH�D$ H��$�   M��M��H�D$(tH�t$ H���i ��t/M9�tNA�9�rKH�t$ �I��M9�t7A�9�r4H���hl ��u�   H�T$pH�L$ L�H��$�   H�
H��8[^�1��ݸ   �֐����UWVSH��8�AL��$�   �yL��L�D$ L�L$(u<I�Z�M��t"H�l$ ��H���i 9���H����H����u�H�D$ H)�H��8[^_]�H�l$ H���Qn 뵐���������������A����������Ð�������������H��XH��$�   L�D$0D�AH�T$@L�L$8D�IH�L$0H�D$@H��$�   �D$    A��A����  H�D$H���  DC�A����n H��$�   H�L$0H�
H��$�   H�L$@H�
H��XÐ�����������H��XH��$�   L�D$0D�AH��H�T$@H��$�   H�L$0L�L$8�D$    D�HA����  H�T$H���  DC�H�T$@�p H��$�   H�L$0H�
H��$�   H�L$@H�
H��XÐSH��0�AL��L�ʉD$ L�D$`D�IH���=o H)�H��0[Ð����A����������Ð�������������H��XH��$�   L�D$0D�AH��H�T$@H��$�   H�L$0L�L$8�D$    D�HA����  H�T$H���  DC�H�T$@�vm H��$�   H�L$0H�
H��$�   H�L$@H�
H��XÐH��XH��$�   L�D$@D�AH��H�T$0H��$�   H�L$@L�L$H�D$    D�HA����  H�T$8���  DC�H�T$0�6o H��$�   H�L$@H�
H��$�   H�L$0H�
H��XÐSH��0�AL��L�ʉD$ L�D$`D�IH����m H)�H��0[Ð���WVSH�� H��H��H��L���c ��tH� H�� [^_��     I��H��H��       �H�� [^_���������������WVSH�� H��H�	��@��H����@ ���u.�z�H�
��H���� ؉�uH@8���H�� [^_�f.�     1�H�AH9Ar�H�H�T$H�PHH�T$H���u�H�    ���@ 1�H�AH9Ar�H�H�T$H�PHH�T$H���u�H�    ��댐���SH�� ���H�ˉ�H�	uH��u	H�� [� H�AH;As	� H�� [�H��PH���u�H�    �А��������SH�� ���H�ˉ�H�	uH��u	H�� [� H�AH;As	� H�� [�H��PH���u�H�    �А��������WVSH�� H��H�	f����H���� ؉�u/f�z�H�
A��H����D ���u6D8���H�� [^_��     H�AH;AsJ� 1�f���u�H�    ���H�AH;As� E1�f���u�H�    A���H�H�T$H�PHH�T$H��H�H�T$H�PHH�T$H말���������SH�� f���H�ˉ�H�	uH��uH�� [�f�H�AH;As� f���u�H�    ��@ H��PH�吐������SH�� f���H�ˉ�H�	uH��uH�� [�f�H�AH;As� f���u�H�    ��@ H��PH�吐�������A����������Ð�������������ATUWVSH��@�A�qH��$�   H��$�   H�|$0�D$,M��H�T$,H��L�D$0L�L$8�=b H�T$0H�D$8H)�H��vkH9�u'�   9���   H���C�H�D$8H)�H��vDH9�tnD�D$,��H���d H�T$0���uŸ   H��$�   H��$�   H�H�H��@[^_]A\�H��$�   H�H��$�   H�1�L9����H��@[^_]A\�@ H��$�   H�H��$�   H��   H��@[�       ^_]A\�f.�     �   �v���������VSH��8H�D$x�q�YH�D$ H�L$ M��M��H��$�   ��H�D$(�a H�L$ ��t(M9���   A�9�rc��L�D$(I)�=��  w`I��w�   H�T$pL�H��$�   H�
H��8[^É�f����D�I��M9�f�H�D$ H�HH�L$ tbA�9�s��   ��     I��v�A��f%�A��
f- $fA��@(��t4fD�H�L$ H�QH�T$ f�AH�D$ I��M9�H�HH�L$ u�1��X���fA��f��fD�H�L$ H�QH�T$ ��ATUWVSH��@H��$�   �AD�aH�l$0L��L�D$0H�T$,H��L�L$8�D$,H�_���_ H��t$D�D$,D��H���kb H����A9���H����u�H�D$0H)�H��@[^_]A\Ð����A����������Ð�������������SH��@H�T$xH��H�T$0H��$�   L��L�D$ D�@H�L$ L�L$(D�HH�T$8H�T$0�c H�L$pH�T$ ��L�D$0H�H��$�   L�uH9ں   E�H��@[Ð����������SH��@H�D$xD�Y�YH�D$0H��$�   L�T$0D��L��L�D$ L�L$(H�D$8�S_ �   ��tL��E��A��H�L$ ��d ��H�D$pH�L$ H�H��$�   H�L$0H���H��@[�SH��0H�T$`H��L��L�D$ L�L$(D�@H�L$ D�H�$g H)�H��0[Ð�����������A����������Ð�������������SH��@H�T$xH��H�T$0H��$�   L��L�D$ D�@H�L$ L�L$(D�HH�T$8H�T$0�Mb H�L$pH�T$ ��L�D$0H�H��$�   L�uH9ں   E�H��@[Ð����������SH��@H�D$xD�Y�YH�D$ H��$�   L�T$ D��L��       �L�D$0L�L$8H�D$(��] �   ��tL��E��A��H�L$0�wc ��H�D$pH�L$0H�H��$�   H�L$ H���H��@[�SH��0H�T$`H��L��L�D$ L�L$(D�@H�L$ D�H��e H)�H��0[Ð����������H�9 Ð��������A����������Ð�������������ATUWVSH��0�AH��$�   H��$�   �qM��L�D$ L�L$(��   H�l$ M9�tAf�H9�t:��H���Q] �����   9���   =��  wH�S�L�d$ H��L�L$(M9�u�1��H��H)�H��u&�   H��$�   L�"H��$�   H�H��0[^_]A\É�f%���
f- $f��@(���҉C�H�S��     H�L$ �a L�d$ L�L$(�;����    L�d$ �   �@ L�d$ �   �u����WVSH��0H�D$x�A�qH�D$ H��$�   M��L��H�D$(tH�L$ �[ ����   H��L)�H��I9���   H�|$ �V�    H����   A�B�� $�����  w[��
A�   �� $��9�rGH���X^ ��tDO��H��L)�H��L9�tVA��� (�����  v��� $��=�  v
9�A�   s��   �f��   H�T$pH�L$ L�H��$�   H�
H��0[^_�1��ܐ������SH��0�AL��L�ʉD$ L�D$`D�IH���Y H)�H��0[Ð����A����������Ð�������������H��XH��$�   L�L$8D�IH��H�T$@H��$�   H�L$0L�D$0�D$     D�@A��H�T$HH�T$@A����` H��$�   H�L$0H�
H��$�   H�L$@H�
H��XÐ��������H��XH��$�   H��H�T$@H��$�   �D$     H�L$0L�D$0D��       @L�L$8D�HH�T$HH�T$@�b H��$�   H�L$0H�
H��$�   H�L$@H�
H��XÐSH��0�AL��L�ʉD$ L�D$`D�IH���MX H)�H��0[Ð����A����������Ð�������������ATUWVSH��0�AH��$�   H��$�   �yL��L�D$ L�L$(��   L�d$ I9�tBf�H9�t;��L���Y �����   9���   =��  wH�Sf�H�t$ H��L�L$(I9�u�1��H��H)�H��u0�   H��$�   H�2H��$�   H�H��0[^_]A\�f.�     ��f%���
f- $f��@(f�Cf�H�S돐H�L$ ��] H�t$ L�L$(�;����    H�t$ �   �@ H�t$ �   �v����WVSH��0H�D$x�A�qH�D$ H��$�   M��L��H�D$(tH�L$ ��W ����   H��L)�H��I9���   H�|$ �W�     H����   A�B�� $�����  w[��
A�   �� $��9�rGH���Z ��tCO�ZH��L)�H��L9�tVA��� (�����  v��� $��=�  v
9�A�   s��   ���   H�T$pH�L$ L�H��$�   H�
H��0[^_�1��ܐ������SH��0�AL��L�ʉD$ L�D$`D�IH����U H)�H��0[Ð���VSH��HH�H�\$ H��H���P L�D$(H��H�T$ �d H�L$ H��H9�t�$� H��H��H[^�H�L$ H��H��H9�t�� H���le��������������SH��0H�H��H�L$(�PH�T$(H��L�B��e H�L$(�������A���~	H��H��0[�H�T$'H���� H��H��0[�H�T$'H��H�D$(H�H��� H����d�������������1�H;Jt��    D9��Ð�       ��������SH��0H�H�@(L��L�J   L9�u%1�H9KtH��0[��    9��H��0[�D  L�L$ A��H��L���ЋT$ H�L$(�������H��D�H�QÐ����UWVSH��(L9�H��H��L��s;H�-C   ���;   H���C�H9�t H�H���H�@ H9�t���H���C�H9�u�H��H��([^_]Ð��H�I0D�� B�AL��E�Ð��������UWVSH��(L9�H��H��L��s;H�-C   ���;   H���C�H9�t H�H���H�@H9�t���H���C�H9�u�H��H��([^_]Ð��H�I0D�� B�AL��E�Ð��������WVSH��   1�H�\$ H�ΈH��H=   u�H�H��  H�~9H�@8H9�u9A�   H��H������F8A�   H��H����
����t�F8H��   [^_�I��H��H��L��$   ���Ð�������UWVSH��H  1�H�\$@H�ΈH��H=   u�H�H�-�  H��9  H�@HH9�u\A�   H��H���q
��Ɔ9  A�   H��H���a
����uH�H�@HH9�u=�D$@�D$?�|$?uƆ9  H��H  [^_]�H�|$ E1�H��H��L��$@  ���H�T$?A�   H��H�T$ L�CH����뮐�������������VSH��8�A8<H��L��t��t+H�H��   H�@8H9�u5I��L��I)��	��H��H��8[^�L�L$(H�T$ �>���L�L$(H�T$ �f�I��H��H��8[^H���VSH��(H�ˉ�����H�H�F   H�@0H9�u��H��([^�@ @��H��H��([^H��SH�� L��L��I)��	��H��H�� [Ð�����Ð������������SH�� H�L$PL��I)�����H��H�� [Ð���Ð�������������       UWVSH��(M9�H��L��s5��L���D  H��H9�vH���H��D��P��t�H��H��([^_]�L����WVSH�� L9�H��L��s$I�@�H)�H��H�tB�H������f�C�H9�u�H��H�� [^_Ð���������������������������WVSH�� L9�H��L��s$I�@�H)�H��H�tB�H���[��f�C�H9�u�H��H�� [^_Ð�����������������0����������UWVSH��(M9�H��L��s5��L���D  H��H9�vH���H��D��P��u�H��H��([^_]�L����f����   v4f�� ��   wWf�� ��   f��@��   H��� �7u���    f����   wDf����   f����   H��� �u��@ f�� ��   f��u^H��� ��t��f�f����   f��u@H��� ��t��@ H��� �t��@ H�M� �t��@ H�1� �t��@ f�� tI1��fD  H�/� �tt��@ H�� �dt��@ H�� �Tt��@ H�� �Dt��@ H�� �4t������AWAVAUATUWVSH��(L9�H��M��M��sUI�@�L���  H)�H���  H��M�tAD  L��1��S ������tf;H��H9�u�fA�<$I��H��M9�u�L��H��([^_]A\A]A^A_Ð��������UWVSH��(H���  ��A��H���  �f�H��H9�t'f�;t��S �������t�   H��([^_]�D  1�H��([^_]Ð����SL9�s&L��E1�H)ӐF�F��Y�   fG�QI��L9�u�L��[Ð������������������Q�   Ð���AUATUWVSH��(�y H��$�   �       I��H��L��D��tjL9�sRI�@�H)�H��L�lB�@ Hc�H��H��A�D�F�I9�t$�f��v��	r�����D�H��H���F�I9�u�H��H��([^_]A\A]� L9�s�I�@�H)�H��L�d���q�����D�H��H���F�L9�u�H��H��([^_]A\A]Ð�������������SH�� f��D����w�y u���rq�����D�H�� [�fD  �DH�� [Ð����H�H��tH��� �   ���� ��H�H�H��Ð�����AWAVAUATUWVSH��8�A H�H�iH��H�)I��H�A    L�h M�u M���c  I�} �  L��1� H��I�|� H������H��H��A������A�tڅ���  ��   H���%z H�~  L�0I�6H�����H��������H+KI��H9��2  H��H���{{ H�H�sH9�H�~�	  H�SH9���  �0=H�H�{�D0 I�$H�@ H�0H���'��H��������H+KI��H9���  H��H���{ I���������   H�H�{H9�L��2  H�SI9���   �8;H�L�{�D8 I�<6H�����I��L��H+CI9��w  H��H���z H�H�{H9�L���   H�SI9���   �8=H�L�{�D8 I�$H�@ H�<0H���S��I��L��H+CI9��  H��H���Ez H��H��0�4���H��H��8[^_]A\A]A^A_� H�D$    E1�E1�H��H����{ H�����H�D$    E1�E1�H��H���{ H��U���L���� ��M��E1�1�H�D$ H����] 놺   ����� �   ����fD  �D$ *   A�   E1�1���d �L��� �       H�D$    E1�E1�H��H���&{ H������   �����H�� ��A H��� �A H��� �A H��� �A H�H��H9�t�� H���lX��������������AVAUATUWVSH��@L�d$?H��H��1�1�M���� H�U H�L�j M�u M����  I�} ��  L��1� H��I�|� H������H��H��A������A�tڅ���  ��   H���e H�> L�(I�u H���O���H��H��I���! H�H�x�H�wH;p��0  H��H���! H�H�P��=H�H�p��@�    �D8 H�E H�@ H�0H�������H��H��I���� �   H�L�p�I�~H;x�w�@���~H��H��� H�H�P��;H�H�x��@�    B�D0 I�|5 H������H��H��I���` H�L�p�I�~H;x�w�@���~H��H���] H�H�P��=H�H�x��@�    B�D0 H�E H�@ H�<0H���*���H��H��I����
 H��H��0�1���H��H��@[^_]A\A]A^Ë@�������������L�������L��H��I��� ��@ L�@�A�   1�H���D$ *   �t �H�H��L��H���� H���V����������WVSH�� L��< I������H��H��H��< �i� H��tH�H��H�� [^_�fD  H;Y ��   H;� �&  H;_ ��  H;� �O  H;� �  H;� ��  H;{ ��  H;� �X  H; �{  H;D �x  H; �  H;J �K  H;] �x  H;P ��  H;3 �t  H;� �C  �(   趍�        1�H��H���y H�s ��FH�9~ H���������   膍 1�H���@    H�3  f�OH�(   H�G    H�G    H���G  H�H�G(    H�G0    H�G8    H�G@    Ƈ�    �#� 1�H���@    H�@! H�{H��H��H�� H�s��FH�~ 1�H�I��H��H�{ 蹍 �3���@ �   �ƌ H���@    H�! H�sH��H���FH��~ H�������    茌 H���@    H�K  H��H��oE H�CH�s��FH��{ H����� �    �F� H���@    H�� H��H��)E H�CH�s��FH�5{ H��l����   �� H���@    H��  H�sH��H���FH�� H��2��� �   �Ƌ H���@    H��  H�sH��H���FH�� H������fD  �p   膋 1ҹ(   H���@    H�� f�W H�G    H�G    H���G" H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Go �� E1�1�H���@    H�Q H�{H��H��H��n# H�s��FH�� 1�H�I��H��H�{ �j� ����D  �p   覊 �(   H���@    H�� H�G    H�G    �G" H��H�G(    H�1�f�G H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Go �'� E1�1�H���@    H�a H�{H��H��H��� H�s��FH�. 1�H�I��H��H�{ �Z� �4���D  �(   �Ɖ 1�H��H�       ��� H�s ��FH��y H�� ������   薉 �(   H���@    H�P H�G    H�G    �G  H��H�G(    H�H�G0    H�G8    H�G@    �GH    Ƈ�    �2� 1�H���@    H�_ H�{H��H��H��L H�s��FH��z 1�H�I��H��H�{ �h� �B����   �و H���@    H�( H�sH��H���FH��{ H������   蟈 H���@    H�^ H�sH��H���FH��| H�������   �e� H���@    H�D H�sH��H���FH�} H�������   �+� �(   H���@    H�U H�G    H�G    �G  H���G"    H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Gz 談 E1�1�H���@    H� H�{H��H��H��' H�s��FH�R 1�H�I��H��H�{ �� ������   �O� �(   H���@    H�i H�G    H�G    �G  H���G"    H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Gz �φ E1�1�H���@    H�) H�{H��H��H���" H�s��FH��} 1�H�I��H��H�{ �� �����H�� �5 H�KH���
  H���-& H���� H���}M��H��H���@ ��H�KH����	  H��� ������H����H�KH����	  H���) ��H�KH���	  H���� �H��H���? H��蠅 H���M��H�KH���|	  H���        �b����m���H�KH���^	  H���! �D����O�����o��������WVSH�� L�r3 I������H��H��H�n3 �)� H��tH�H��H�� [^_�fD  H;� ��   H;\ �&  H;� ��  H;� �O  H;� �  H;� ��  H;� ��  H;. �X  H;Q �{  H; �x  H;W �  H;j �K  H;} �x  H;� ��  H;� �t  H;� �C  �(   �v� 1�H��H����� H�s ��FH�9u H���������   �F� 1�H���@    H�� f�OH�(   H�G    H�G    H���G  H�H�G(    H�G0    H�G8    H�G@    Ƈ�    �� 1�H���@    H�p H�{H��H��H��� H�s��FH�u 1�H�I��H��H�{ 詂 �3���@ �   膃 H���@    H�5 H�sH��H���FH�v H�������    �L� H���@    H�� H��H��/< H�CH�s��FH��r H����� �    �� H���@    H�u H��H���; H�CH�s��FH�5r H��l����   �Â H���@    H�� H�sH��H���FH��v H��2��� �   膂 H���@    H�u H�sH��H���FH�w H������fD  �p   �F� 1ҹ(   H���@    H�N f�W H�G    H�G    H���G" H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �       �Go �ǁ E1�1�H���@    H� H�{H��H��H���A H�s��FH�x 1�H�I��H��H�{ �ڋ ����D  �p   �f� �(   H���@    H�` H�G    H�G    �G" H��H�G(    H�1�f�G H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Go �� E1�1�H���@    H� H�{H��H��H��N= H�s��FH�^v 1�H�I��H��H�{ �ʆ �4���D  �(   膀 1�H��H���)� H�s ��FH��p H�� ������   �V� �(   H���@    H� H�G    H�G    �G  H��H�G(    H�H�G0    H�G8    H�G@    �GH    Ƈ�    �� 1�H���@    H�� H�{H��H��H��� H�s��FH��q 1�H�I��H��H�{ ��� �B����   � H���@    H�X H�sH��H���FH��r H������   �_ H���@    H�> H�sH��H���FH��s H�������   �% H���@    H�$ H�sH��H���FH�t H�������   ��~ �(   H���@    H� H�G    H�G    �G  H���G"    H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Gz �k~ E1�1�H���@    H�� H�{H��H��H��"F H�s��FH��v 1�H�I��H��H�{ �� ������   �~ �(   H���@    H�) H�G    H�G    �G  H���G"    H��       H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Gz �} E1�1�H���@    H�� H�{H��H��H��vA H�s��FH��t 1�H�I��H��H�{ �ҋ �����H��� �q, H�KH����   H���D H����| H���=D��H��H����6 ��H�KH���   H����� ������H����H�KH���   H���-H ��H�KH���m   H���U� �H��H���x6 H���`| H����C��H�KH���<   H���< �b����m���H�KH���   H���&@ �D����O�����o����������it	��     H�H�`���������UWVSH��xH�H��H�H��H9���   H�x H�H����   H�j H�U H��t{�������urH� tvH�|$PH��H���f���H�t$0H��H���V���L�D$81�L;D$XH�\$0tXH��H9�tH�وD$/�^{ �D$/H�L$PH��H9�t�D$/�B{ �D$/�1�H��x[^_]�H�} u��   H��x[^_]�M���   t�H�T$PH���|��������H�L$PH��H��H��H9�t��z H��H��H��u
��} H�����9B�����������H�y  H�H�@PH9�uH�A�@`�D  H���������������H�Y  H�H�@HH9�uH�A�@\�D  H���������������VSH��(H�H�@(H��H�9  H9�uDH�BI������H�p(H�CH�H��tH���!���L�E1�H��H���K H��H��([^�D  H����H��H��([^ÐVSH��(I������H�BH�pH�AH��H�H��tH�������L�E1�H��H���J H��H��([^Ð��������       H��  H�H�@@H9�uH�A�@X�D  H���������������H��  H�H�@H9�uH�A�@!�@ H���������������H�A�@`Ð�������H�A�@\Ð�������VSH��(H�H�@8H��H�i  H9�uDH�BI������H�pHH�CH�H��tH�������L�E1�H��H����I H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�I  H9�uDH�BI������H�p8H�CH�H��tH���q���L�E1�H��H���_I H��H��([^�D  H����H��H��([^ÐH�9  H�H�@H9�uH�A�@"�@ H���������������VSH��(I������H�BH�p(H�AH��H�H��tH�������L�E1�H��H����H H��H��([^Ð�������H�A�@XÐ�������H�A�@!Ð������VSH��(I������H�BH�pHH�AH��H�H��tH���t���L�E1�H��H���bH H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH���$���L�E1�H��H���H H��H��([^Ð�������H�A�@"Ð������VSH��(H�H�@ H��H�����H9�uDH�BI������H�pH�CH�H��tH������L�E1�H��H���G H��H��([^�D  H����H��H��([^ÐH�y  H�H�@PH9�uH�A�@`�D  H���������������H�Y  H�H�@HH9�uH�A�@\�D  H���������������VSH��(H�H�@(H��H�9  H9�uDH�BI������H�p(H�CH�H��tH�������L�E1�H��H����F H��H��([^�D  H����H��H��([^ÐVSH��(IǤ       �����H�BH�pH�AH��H�H��tH������L�E1�H��H���rF H��H��([^Ð�������H��  H�H�@@H9�uH�A�@X�D  H���������������H��  H�H�@H9�uH�A�@!�@ H���������������H�A�@`Ð�������H�A�@\Ð�������VSH��(H�H�@8H��H�i  H9�uDH�BI������H�pHH�CH�H��tH������L�E1�H��H���E H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�I  H9�uDH�BI������H�p8H�CH�H��tH���1���L�E1�H��H���E H��H��([^�D  H����H��H��([^ÐH�9  H�H�@H9�uH�A�@"�@ H���������������VSH��(I������H�BH�p(H�AH��H�H��tH������L�E1�H��H���D H��H��([^Ð�������H�A�@XÐ�������H�A�@!Ð������VSH��(I������H�BH�pHH�AH��H�H��tH���4���L�E1�H��H���"D H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH�������L�E1�H��H����C H��H��([^Ð�������H�A�@"Ð������VSH��(H�H�@ H��H�����H9�uDH�BI������H�pH�CH�H��tH���q���L�E1�H��H���_C H��H��([^�D  H����H��H��([^ÐH�y  H�H�@PH9�uH�A�@`�D  H���������������H�Y  H�H�@HH9�uH�A�@\�D  H���������������VSH��(H�H�@(H��H�9  H9�uDH�BI������H�p(H�CH�       �H��tH���I���L�FE1�H��H����j H��H��([^�D  H����H��H��([^ÐVSH��(I������H�BH�pH�AH��H�H��tH���D���L�E1�H��H���2B H��H��([^Ð�������H��  H�H�@@H9�uH�A�@X�D  H���������������H��  H�H�@H9�uH�A�@"�@ H���������������H�A�@`Ð�������H�A�@\Ð�������VSH��(H�H�@8H��H�i  H9�uDH�BI������H�pHH�CH�H��tH���	���L�FE1�H��H���i H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�I  H9�uDH�BI������H�p8H�CH�H��tH������L�FE1�H��H���/i H��H��([^�D  H����H��H��([^ÐH�9  H�H�@H9�uH�A�@$�@ H���������������VSH��(I������H�BH�p(H�AH��H�H��tH������L�FE1�H��H���h H��H��([^Ð�������H�A�@XÐ�������H�A�@"Ð������VSH��(I������H�BH�pHH�AH��H�H��tH������L�FE1�H��H���2h H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH���L���L�FE1�H��H����g H��H��([^Ð�������H�A�@$Ð������VSH��(H�H�@ H��H�����H9�uDH�BI������H�pH�CH�H��tH���1���L�E1�H��H���? H��H��([^�D  H����H��H��([^ÐH�y  H�H�@PH9�uH�A�@`�D  H���������������H�Y  H�H�@HH9�uH�A��       @\�D  H���������������VSH��(H�H�@(H��H�9  H9�uDH�BI������H�p(H�CH�H��tH���	���L�FE1�H��H���f H��H��([^�D  H����H��H��([^ÐVSH��(I������H�BH�pH�AH��H�H��tH������L�E1�H��H����= H��H��([^Ð�������H��  H�H�@@H9�uH�A�@X�D  H���������������H��  H�H�@H9�uH�A�@"�@ H���������������H�A�@`Ð�������H�A�@\Ð�������VSH��(H�H�@8H��H�i  H9�uDH�BI������H�pHH�CH�H��tH�������L�FE1�H��H���_e H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�I  H9�uDH�BI������H�p8H�CH�H��tH���Y���L�FE1�H��H����d H��H��([^�D  H����H��H��([^ÐH�9  H�H�@H9�uH�A�@$�@ H���������������VSH��(I������H�BH�p(H�AH��H�H��tH�������L�FE1�H��H���bd H��H��([^Ð�������H�A�@XÐ�������H�A�@"Ð������VSH��(I������H�BH�pHH�AH��H�H��tH���\���L�FE1�H��H����c H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH������L�FE1�H��H���c H��H��([^Ð�������H�A�@$Ð������VSH��(H�H�@ H��H�����H9�uDH�BI������H�pH�CH�H��tH�������L�E1�H��H����: H��H��([^�D  H����H��H��([^Ð�       �   L�I9�w
LAL9���Ð�������H�AH9��Ð����WVSH�� H��H��H��L���x���I��H��H��I��H�� [^_�    UWVSH��(H�AH��H��L��tIM��tDH��L��H�)L9�HF���H��H���t�T I��H������H��t�H��H��([^_]�D  H������H��H��([^_]Ð������������L�JH��t�������H������L�IM��tL�H�	I9�IF� :t
H��H���u��H�AÐ����������WVSH�� H��H��H��L���x���I��H��H��I��H�� [^_�    ATUWVSH�� M��H��L��L��tHH�yI9�s?L�!�f.�     H��H9�t'A�I��H������H��t�H��H�� [^_]A\�@ H������H�� [^_]A\Ð�������������L�JH��t����������(  ��������H��Ð�����������H��(I��������L�H+QL9�rH��(�L��� ���������H��Ð�����������WVSH�� H��H��H��L���X���I��H��H��I��H�� [^_�    UWVSH��(H������H�AH��H��L��t1H�H�)L9�IG�H��t�T I��H������H��t
H��H���u�H��H��([^_]Ð����L�JH���������H������L�IM��tL�H�	L9�IG���H��H���t8t��WVSH�� H��H��H��L������I��H��H��I��H�� [^_�    ATUWVSH�� H�yI9�H��L��L��sDM��L�!u�(f.�     H��H9�t'A�I��H������H��u�H��H�� [^_]A\�@ H������H�� [^_]A\Ð�������������L�JH��t�������H������L�IM9�A��s#H�B:�        t
�"f�F8 uI��M9�u�H�������f�     L��Ð�����������H��(L�AL9�sH�H�H��(�H�Q� �, ������������H�AHÐ�������H�AH�H�D�Ð��H�AHÐ�������SH�� H�YI9�H��L��w:L)�L9�IG�H��tHH��tI��H���i���H��H�� [���H��H�� [�H��� I��I��H��� � ���������H�Ð�����������WVSH�� H��H��H��L������I��H��H��I��H�� [^_�    AVAUATUWVSH�� M��H��L��H�Q��   L9�H������vgH�)H�| L)�J�L I9�wRA�   M)�L�I��tAD�.D������H��I��t&I��H��H��������tGI�NI��I)�L9�wM�u�H������H�� [^_]A\A]A^�L9�H������IC�H�� [^_]A\A]A^�L��H)��̐�������L�JH��$�������VSH��(H������H�AI9�s"H�1L)���J�I�������H��H)�H��HE�H��H��([^Ð�������������H�H��H�Ð�����H�AÐ����������H�Ð�����������H�Ð�����������H�H��H�Ð�����H�y ��Ð������H�Ð�����������WVSH�� H��H��H��L�������I��H��H��I��H�� [^_�    UWVSH��(H������H�AI9�H��L��w:L)�L��H�)L9�HF�H��t%H�L I��H���������tH�C�H��tH��H��u�H��H��([^_]�H�������됐�L�JH���������H������L�IM��tL�H�	L9�IG� 8t
H��H���u��H�Ð�����������H�AÐ����������L�BLH��L�Ð��       SH�� H�BI9�H��w9H�AH�H�JH�I9�w<J� L)�L9�IG�E1�L�
H���2 H��H�� [�H�ó I��H�� �0 H��� I��H�� � ����������H�Ð�����������UWVSH��(H�YH��H��H���&���I��H9�H��LF�M��tH�H��������uH)����H������@H��   �M�H��([^_]Ð�������������VSH��(H�YH�rI��H9�LF�M��tH�H�	� �����uH)����H������@H��   �M�H��([^Ð��������������ATUWVSH�� H�YH9�H��H��M��w`H)�L��L9�IG��B���H9�I��H��LF�M��tHu L��H��������uH)�����H������@H��   �M�H�� [^_]A\�H��� I��I��H��� � �����������VSH��(H�YH�t$`H9�wPH)�L9�IG�I��H9�LF�M��tHH��L��������uH)����H������@H��   �M�H��([^�H�� I��I��H�.� � ���VSH��(H�YH9�wTH)�I�qL9�IG�H9�I��LF�M��tHH��I�������uH)����H������@H��   �M�H��([^�H��� I��I��H��� � ����VSH��(H�YL�T$hH��H�T$`H9�wcI�qH9�wsH)�L9�IG�H)�L9�IG�I��H9�LF�M��tHIH���������uH)����H������@H��   �M�H��([^�H� � I��I��H�� �� H�ٮ I��I��H��� �� ���������������L�BLH��L�Ð�H��(L�IH��L��L9�wH��(�H��� I��� ��       ��������H�AH)�L9�IG�ÐH�AH9tH�A�f��   Ð���������H��������Ð����H�H�Ð���������   L�I9�wH�AI�@H9���Ð���H�AH9��Ð����WVSH�� H��H��H��L�������I��H��H��I��H�� [^_�    H�AH��tBM��t=H��L�L9�IG�@ H��E�CtH��M��fD;tH��I��u�H��H���u��H������Ð������������L�JH���������H������L�IM��t L�H�	I9�IF� f;At
H��H���u�Ð��������������H�AÐ����������WVSH�� H��H��H��L�������H��t<H�WH9�s3L��    H��E�[tH��I��fD;tH��I��u�H��H9�u�H������H��H�� [^_Ð����VSM��tBH�YI9�s9H�1L��f.�     H��D�FtH��M��fD;tH��I��u�H��H9�u�H������[^Ð������������VSH�rL�H��t;L�YM9�s2H�L�� M��D�CtL��H��fD;
tH��H��u�H��L9�u�H������[^Ð������������H������L�IM9�s)L�L��L)�O�BM��tfA;tI��H��u�H�������fD  M)�L��H��Ð�����H��Ð�����������H��(I��������?L�H+QL9�rH��(�L���9 ���������H��Ð�����������WVSH�� H��H��H��L��� ���I��H��H��I��H�� [^_�    H������L�QM��t2L�L�L9�IG�M��t H��E�CtH��M��fD;tH��I��u��H��H���u�Ð�L�JH���������H������L�IM��t L�H�	L9�IG����       H��H���tf9At�Ð��������������WVSH�� H��H��H��L���P���H�WH9�sOL�H��I�Xt#H��D�tH��I��@ fD9tH��I��u�H��H�� [^_�D  H��H9�tE�X��H�������א������SH�AI9�sFH�M��J�CtH��D�tH��M��fD9tH��I��u�L��[�fD  I��L9�tF�C��I�������ܐ������SL�QH�BM9�sGL�H��K�Ct&H�D�	H��tH��H��@ fD9
tH��H��u�L��[�I��M9�tG�C��I�������␐H������L�IM9�A��s$H�fB;@t
�!�fF9@uI��M9�u�H��������     L��Ð�����������H��(L�AL9�sH�H�PH��(�H�p� �� �����������H�QH�H�PÐ���H�QH�H�DP�Ð��H�QH�H�PÐ���SH�� H�YI9�I��L��wAL)�L9�IG�H��tH�H��J�JtL�L������H��H�� [��fA�H��H�� [�H��� I��I��H��� �" ��H�Ð�����������WVSH�� H��H��H��L�������I��H��H��I��H�� [^_�    WVSL�YM����   M9�H������vKH�1L��L)�I9�N�Fw9�   L)�M��H�t!H��t�
J�<^M�Y��fA;
tI��H��u�H������[^_�D  L9�tM1�L9�tFE�DBH��fD;Bt�I��H��L)�H��I9�w�H�M��t�H��u��f�M9�H������IC�[^_�L��H)�H��뚐��L�JH��$�������H������L�IM9�s)L�L��L)�O�BM��tfA9tI��H��u�H�������fD  M)�L��H��Ð�����H�H��H��       Ð�����H�AÐ����������H�Ð�����������H�Ð�����������H�H��H�Ð�����H�y ��Ð������H�Ð�����������WVSH�� H��H��H��L������I��H��H��I��H�� [^_�    H������L�QM9�wWH�	M�Y�M)�L��M9�IF�L�AM��t:I9�t5M��A��H����A8�u,�
fA9u#1��E�THH��fD;JuI9�u���     H�H�I��H��tH���H������Ð�����L�JH��d�������H������L�IM��t L�H�	L9�IG� f9At
H��H���u�Ð��������������H�Ð�����������H�AÐ����������H��H�JH�H�JH�Ð�������������SH�� H��H�JI9�w0H�CL)�H�H�L9�IG�E1�J�@L�JH���HM H��H�� [�H��� I��H�� �
 ���������H�Ð�����������WVSH�� H�YH��H��H���O���H��H9�HF�H��tXL�L9�tPM��A��H����A8�tH�������H�� [^_�f.�     1��<NfA9<HuCH��H9�u�f.�     H)ø���H������@H��   �M�H�� [^_�f.�     ���H�� [^_Ð��H�AL�BI��I9�MF�M��tIL�H�	I9�t>H��A��M����A8�tI��������1�E�RfD9Qu3H��L9�u��     L)�H�¸���H�����̍@H��   �M�����Ð�������UWVSH��(H�YH9�H��H��L����   H)�L��L9�IG������H9�H��HF�H��tQH�U L�zI9�tDM��A��H����A8�tH�������H��([^_]�1��<VfA9<Pu@�       H��H9�u��    H)ø���H������@H��   �M�H��([^_]�f�     ���H��([^_]�H�å I��I��H�� �I ���������H��(H�AL�T$PH9���   H)�M��L9�LF�M9�MF�M��tQH�H�PL9�tEH����M����8�tI�������H��(�@ 1�A�Af9Bu7H��L9�u�f.�     M)и���I������@I��   �AM�H��(����H��(�H�� I��I��H�� �y ���������H��(H�AH9���   H)�M�QL9�LF�M9�M��MF�M��tRH�M�	H�PL9�tCH����M����8�tI�������H��(�f�1�A�Af9Bu7H��I9�u�f.�     M)и���I������@I��   �AM�H��(����H��(�H�#� I��I��H�D� � ���������SH�� L�QL�\$PH�\$XL9���   I�AI9���   I)�M9�MF�L)�H9�HG�M��L9�LF�M��tTM�	H�	O�YH�QI9�tAH��A��M����A8�tI�������H�� [�1�A�Qf9Qu5H��L9�u��    I)�����I������@I��   �AM�H�� [����H�� [�H�1� I��M��H�R� � H�F� I��M��H�� � ��������������H��H�JH�H�JH�Ð�������������H��(L�IH��L��L9�wH��(�H��� I���I ���������H�AH)�L9�IG�ÐH�AH9tH�A�f��   Ð���������H��������?Ð����H�H�PÐ�������H��(H��L���9�������������	�H��(Ð������������AWAVAUAT�       UWVSH��hL�t$ L��I��I�FE1�L��H�D$ L�|$@�� I�GE1�H��L��$�   L��H�D$@� H�\$ H�l$(H�t$@L�d$HH�I��3�H��舼��H��H��}���H�H9�uI9�t&H9�t[I9�tfH��H��I��H��L��� �������t�H�L$@I��L9�t�7M H�L$ I��L9�t�$M ��H��h[^_]A\A]A^A_Ð������f�     �   �H�L$ I��H��L9�t��L H���K�������������H��L��M��骻����AWAVAUATUWVSH��xH�AL��L���A H�H��I��E1�H�A    H�L$PI��H��H�D$@H�AH�L$HH�D$P�k H�|$PH)�H�D$XH�H��H�H�D$8�kL I��������H���B�  H�L�kB�D  I��I��H��L���I���H9�w(H�pH����K H��� L I��I��H��L��H������L��H+SH9���   I��H��H����3 H���ƺ��H�H9|$8t\H��L�cH�H9D$@M�l$t5H�SI9��\���H�D$    E1�E1�L��H���N5 H��:���fD  �   ��f�     H���HK H�D$HH�L$PH��H9�t�@K H��H��x[^_]A\A]A^A_�H��� �� H���XM �T H���H���fO H�D$HH�L$PH��H9�t��J H�H9L$@t��J H���G��H����H���
M H���J �L�9   H�H�@ L9�u�(   �     H���������������H�H�`���������1�L9�sf�     �
��H���I9�u�Ð�������������SH�� H�H���PH��H�� [Ð��������H��(H��L���ٸ������������	�H��(Ð�������������       AWAVAUATUWVSH��hL�t$ L��I��I�FE1�L��H�D$ L�|$@�C I�GE1�H��L��$�   L��H�D$@��B H�D$(H�\$ H�t$@H�,CH�D$HL�$F�4H���/���H��H�C�#���H9�H�4FuI9�t&H9�tZI9�tcH��H��I��H��L����������t�H�L$@I��L9�t�4I H�L$ I��L9�t�!I ��H��h[^_]A\A]A^A_ÿ�������    �   �H�L$ I��H��L9�t��H H���K�������������H��L��M���b�����AWAVAUATUWVSH��xH�AL��E1�H�A    L��H�H��I��fD�AH�L$PE1�I��H�D$@H�AH��H�L$HH�D$P�A H�\$PH)�H�D$XH�CH�D$8H��������?H9���  H�?�UH I��������?H���fD  1�1�fB�`L�nfB�L`I��I��H��L���,���H9�w<H�xH����G H��������?H9���   H�?��G I��I��H��L��H�������L��H+VH9���   I��H��H���Y H���=���H�CH9\$8tZH��L�fH�H9D$@M�l$t3H�VI9��F���H�D$    E1�E1�L��H���Z H��$���@ �   ��f�     H���G H�D$HH�L$PH��H9�t�G H��H��x[^_]A\A]A^A_�H�%� �� H���(I ��O �P H���6K H�D$HH�L$PH��H9�t�F H�H9L$@t�F H�����H�����]P H����H����H H���xF 랐�����L�9   H�H�@ L9�u�(   �     H���������������H�H�`���������1�L9�sf�     �
��H���I9�w�Ð�������������SH�� H��       H���PH��H�� [Ð��������H�Ð�����������H�QH��H�A    H��A Ð��������SH��0H�H��H�L$hH�L$(�L$`�L$ H���PH��H��0[Ð���L��   H�H�@L9�u1��f.�     H���������������L�y   H�H�@L9�u1��f.�     H���������������L�Y   H�H�@ L9�u�H�����������SH�� E1�H�D$XH�QH��H�H�L�@I�� H��H�� [Ð1�Ð������������Ð��������������H�Ð�����������H�QH��H�A    H�1�f�QÐ������SH��0H�H��H�L$hH�L$(�L$`�L$ H���PH��H��0[Ð���L��   H�H�@L9�u1��f.�     H���������������L�y   H�H�@L9�u1��f.�     H���������������L�Y   H�H�@ L9�u�H�����������SH�� E1�H�D$XH�QH��H�H�H�@L�B�= H��H�� [�1�Ð������������Ð��������������VSH��(I������H�BH�pH�AH��H�H��tH���d���L�E1�H��H���R H��H��([^Ð�������VSH��(I������H�BH�p(H�AH��H�H��tH������L�E1�H��H��� H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH���ı��L�E1�H��H��� H��H��([^Ð�������H�Y   H�H�@H9�uH�A�@H�@ H���������������H�9   H�H�@H9�uH�A�@I�@ H���������������H�A�@HÐ������H�A�@IÐ������VSH��(H�H�@ H�˱       H�y���H9�uDH�BI������H�pH�CH�H��tH������L�E1�H��H���� H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@(H��H�Y���H9�uDH�BI������H�p(H�CH�H��tH���q���L�E1�H��H���_ H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�9���H9�uDH�BI������H�p8H�CH�H��tH������L�E1�H��H���� H��H��([^�D  H����H��H��([^ÐVSH��(I������H�BH�pH�AH��H�H��tH��褯��L�E1�H��H��� H��H��([^Ð�������VSH��(I������H�BH�p(H�AH��H�H��tH�������L�FE1�H��H���9 H��H��([^Ð�������VSH��(I������H�BH�p8H�AH��H�H��tH��謮��L�FE1�H��H���B9 H��H��([^Ð�������H�Y   H�H�@H9�uH�A�@H�@ H���������������H�9   H�H�@H9�uH�A�@J�@ H���������������H�A�@HÐ������H�A�@JÐ������VSH��(H�H�@ H��H�y���H9�uDH�BI������H�pH�CH�H��tH���!���L�E1�H��H��� H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@(H��H�Y���H9�uDH�BI������H�p(H�CH�H��tH���Y���L�FE1�H��H����7 H��H��([^�D  H����H��H��([^ÐVSH��(H�H�@0H��H�9���H9�uDH�BI������H�p8H�CH�H��tH������L�FE1�H��H���7 H��H��([^�D  H����H�ز       H��([^ÐH��  H�H�@H9�u1��f.�     H���������������AWAVAUATUWVSH��xH��$�   M�8I�XI�9I��I��M�aH���   H��$�   � L��L�|$PH�@H�L$`H�\$XL�L$@H�|$@L�D$PL�d$HH�@H�t$ H�l$(H�D$8H��$�   H�D$0�  �D$hH�    ����L�|$`H!�H	Ã��@��M����@ �A��uSA�����H��t��u$@8�u�M L��M�>I�^H��x[^_]A\A]A^A_�1�H�WH9Wr�H�H���PH������f�1�I�GI9Gr�I�L���PH����    AD�LD�놐��������AWAVAUATUWVSH��xH��$�   M�8I�XI�9I��I��M�aH���   H��$�   �p L��L�|$PH�@H�L$`H�\$XL�L$@H�|$@L�D$PL�d$HH�@ H�t$ H�l$(H�D$8H��$�   H�D$0��  �D$hH�    ����L�|$`H!�H	Ã��@��M����@ �A��uSA�����H��t��u$@8�u�M L��M�>I�^H��x[^_]A\A]A^A_�1�H�WH9Wr�H�H���PH������f�1�I�GI9Gr�I�L���PH����    AD�LD�놐��������AWAVAUATUWVSH��   I�0I�XM�)M�qH��$�   H��H�D$8   L��$  H�D$HH��$  H��$�   �D$0'  L�L$`�D$(    L�D$pH�t$pH�D$@H��$�   H�D$ H�\$xǄ$�       L�l$`L�t$h��  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   D��$�   E�HdE��A������L��$   AH�A�H���@��H����@ �A���|   A�����M��t��u,@8�uA�$H��H�U H�]H�Ĩ   �       [^_]A\A]A^A_� 1�I�uI9ur�I�E H�T$XL���PHH�T$X�������     A�$�q���fD  1�H�FH9F�t���H�H���PH�    ���AD�HE��V�����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[Ð1�Ð������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[ÐAWAVAUATUWVSH��H�
   I�@I�yI�M�9H�D$0A��H��$�   H��$�   H���   �Y
 H��$�   I��tH��$�   ��  �   E�A��1�H����E1�A�����H�D$(A�����H��@��@ ��(  ��A�����M��t����   1�L;�$�   ��  @����  H��t���  D��A��Hc�A��>9  ��u&I�H�@@H;D$(��   ��*�&  A��>9  �ʍA�<	�  �D� �lAЉ���;�$�   ��   �;�$�   ��   ��A��H�C����H;C�  H��H�CI��A����������     I�GI9G�&���I�D�T$<L���T$8�PH�T$8A����̃��D�T$<�������E1������H�CH9C��   1�������    H�CH;C�  �8��������     D�T$8��A�*   L����D�T$8A����̉�*������    H��$�   ueI��u_��dH��$�   �(H�    ����H#D$0I	�H��$�   H�L�`H��H[^_]A\A]A^A_�H�D�T$8H���PPD�T$8A����������f�H��$�   �       �� L;�$�   t��q����H�H��D�T$<�T$8�PH�    �T$8A����̃���    D�T$<E�HD�����D  H�D�T$8H���PHA�����D�T$8���t
����������   �����1������������AWAVAUATUWVSH��  L��$�  I�0I�XI�9I��I��M�aI���   H��$�  �] H��$�   Ǆ$�       H�@L�L$`L�D$pH���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$�   H���   H���   H�t$pH�\$xH��$   L��H��$  H��$�   H�|$`H�D$@H��$�   H�D$(H��$�   H�D$ L�l$8H�D$0   L�d$h��  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   H��$�  D��$�   D�A���A��H����D �A��u|A�����H��t��u,A8�u�M L��I�I�^H��  [^_]A\A]A^A_�D  1�H�wH9wr�H�H�T$XH���PHH�T$X������f�     �M �v����    E1�H�FH9F�s���H�H���PH�    ���ED�HE��U����UAWAVAUATWVSH��hH��$�   H�EhH�]`�Ao �Ao	H�M0L�mXH���   )E�)M�� I��H��   H����6���H�U�H)�H�E�H�U�H�E�H�t$ H���v�����t$H�Ep�H�E0foU�H�e�[^_A\A]A^A_]ËU�H�M�����H�ۉ�t�E1�E1�� I�L���P@8�tI��L9�tK�D� �@�       8�u�F�4�I��I��L9�u�E1�I����   HcA�   I�L� �����H���     Jc�I�L� ����H9�HG�I��M9�w�H�M�H�AH;A��  H��H�AI���E�����I9�����H�Mп   H��t1�H�AH9A��  �}��H�M���H��A��A ��-  @8������1��I��B��I9�A�v3L�<�H�M�IcH��I�D� B�0�E�t	�����   8�u�H��I9�w�I������I���u���H�M�I����X Hc�E�����M�l� ��L������I9�H���.  A������4@8��2���H�M�H�AH;A�   H��H�AI��D�}�I9���   H�U�H�M��l����������H�M�C�t5 �E�H��t����u�H�AH;A��   @:0t������D  H�AH;AsG� ����1�H�AH9A�����H�D�U��U��PH�U����D�U������H�E�    D������H��PH��������H�E�    ���������H��PP����H��PH����>���H�E�    �   �,���H��PP���������H�EP�8����H��PH��������H�E�    ��������������AWAVAUATUWVSH��h  L��$�  I�0I�XI�9I��I��M�aI���   H��$�  �=  H��$�   H�@L�L$`L�D$pH��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$�   H��P  H��$�   H��X  H��$�   H��`  H��$�   H��h  H��$�   H��p  H��$�   H��x  H��$�   H���  H��$�   H���   H��$   H���   H��$  H���   H��$�         H���   H��$  H���   Ǆ$�       H��$   H���   H��$(  H���   H��$0  H��   H��$8  H��  H��$@  H��  H��$H  H��  H��   L�l$8H�D$0   H�t$pH��$P  L��H��$X  H��$�   H�D$@H��$�   H�D$(H��$�   H�D$ H�\$xH�|$`L�d$h�  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   H��$�  D��$�   D�A���A��H����D �A��uwA�����H��t��u'A8�u�M L��I�I�^H��h  [^_]A\A]A^A_�1�H�wH9wr�H�H�T$XH���PHH�T$X������f�     �M �{����    E1�H�FH9F�x���H�H���PH�    ���ED�HE��Z����AWAVAUATUWVSH��H  L�=ƒ��1�H��$�  H��$�  �Ao�AoH���   H��$�  H��H��$�  )�$�   )�$�   ��� H��H�D$X�� H��I���Ӛ����$�   Ǆ$�       H��$�   H�ƃ��@��H����@ �A���}  ��$�   �H��$�   ��H��t����   1�H9���$�   ��  @����  ����  L�$;E�4$H�oC��59  L����u#I�U L�J@M9���  ����   C��59  ��%��   D�$+C��%9  L����u#I�U L�J@M9���  ���  C��%9  ��Ǆ$�       ��E��   ��O��   ��A��8��  H�=�s ��Hc�H���H�AH9A����H��PH�������HǄ$�       �������H��$�   A�<$��$�   H��t	�����   @8��1  ��       �$�   ��$�   H���t���f.�     1�H�AH9A�s���H��PH����d���HǄ$�       D���P���H�o�|;A��=9  H��������I�U L�J@M9��?  ����   A��=9  ��������     ��uH9�tH��$�  �H��$�  fo�$�    H��H  [^_]A\A]A^A_�@ A��E1�L��A���"���H�AH;A�  @:8����������H��H�AǄ$�   ����H�������\���f�H�AH;Ar�H��PPH��$�   ��fD  E1�A��L��A�ф��������$�   ��$�   H��$�   @ H�}�����    H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(   H��$�  H��$�   H�D$ L��$�   L��$�   �Y���D��$�   H��$�   ��$�   E��H��$�   ��$�   �:�����$�   H��$�  �G�#��� H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   L��$�   �D$0;   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ����D��$�   H��$�   ��$�   E��H��$�   ��$�   �j�����$�   H��$�  �G�S��� H��$�   L��L�p I��I�P�肌��H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�    H��$�  L��$�   H��$�  L��$�   H�D$0H��$�   H�D$(H��$�  H�D$ �,���H��$�   ��$�   H��$�   ��$�   ����f�     H��$�   �       H��$�  H�D$8   H�D$HH��$�  H��$�   L��$�   �D$0<   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �����D��$�   H��$�   ��$�   E��H��$�   ��$�   �������$�   H��$�  ������@ H��$�   L��L��n I��I�P�����H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�   �n���H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@ H�D$8�-�����$�   H��$�   H���fx��I�U0���B�����H��$�  L��$�   H�D$0   H��$�  L��$�   L�t$@fo�$�   H��$�   L�d$ fo�$�   L��$�   H�L$pH�D$8H�߰ L��$�   )�$�   )�$�   L�L$`H�D$(L�D$h�#���H��$�   H��$�   H��H��$�   ��$�   ��$�   ��v����$�   ���*�����$�   �$�   ����H���jw��A�}8 A���R  A�EfA8�t*��$�   H���Cw��A�}8 ���  A�Ed@8������H��$�  L�t$HH�|$p�D$0   fo�$�   �D$(    L�L$`L�d$ L�D$h)�$�   H��$�  H�D$@H��fo�$�   H�D$8   )�$�   �W���H��$�   L�t$HH��H��$�  L�d$ L�L$`H�D$8   L�D$h�D$0;   H��$�   ��$�   fo�$�   �D$(    )�$�   ��$�   H��$�  fo�$�   )�$�   H�D$@�����H��$�   ��$�   H��$�   ��$�   ����f.�     ��$�   H��$�   ��u����A��=9  �       ��u#I�M ��L�I@M9��e
  ���=
  A��=9  ��	H��$�   ��	  ��I H��$�   �����Ǆ$�   �����6���fD  H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@����@ H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   )�$�   )�$�   H��$  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ������$�   H��$�   ��$�   ��H��$�   ��$�   �������$�   H��$�  �G����fD  H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   H��$  H��   H��$  H��  H��$   H��  H��$(  H��  H��$0  H��   )�$�   )�$�   H��$8  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ����D��$�   H��$�   ��$�   E��H��$�   ��$�   �@�����$�   H��$�  �G�)���f�     H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0'  L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ������       �$�   H��$�   ��$�   ��H��$�   ��$�   �l���D��$�   H��$�  E�HdE��A������AH��G�B���f�H��$�   L��L��f I��I�P��r���H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�   �����H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(    �����H�D$XH��$�   fo�$�   fo�$�   H�@H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$   H���   H��$  H���   )�$�   )�$�   H��$  ����f.�     H�D$XH��$�   fo�$�   fo�$�   H�@H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$   H��P  H��$  H��X  H��$  H��`  H��$  H��h  H��$   H��p  H��$(  H��x  H��$0  H���  )�$�   )�$�   H��$8  �;���@ H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@0����@ H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �)���D��$�   H��$�   ��$�   E��H��$�   ��$�   �
�����$�   H��$�  �G����� ��$�   H��$�   �,n��I�U0���B �  H��$�   �D$0   fo�$�   H�D$HH��$�  H��$��          fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(
   H��$�  H��$�   H�D$ L��$�   L��$�   �4���H��$�   ��$�   H��$�   ��$�   ��H��$�   ��$�   ��$�   ��������� H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �i���D��$�   H��$�   ��$�   E��H��$�   ��$�   �J�����$�   H��$�  ���G�0�����$�   H��$�   �ll����A��=9  ��u#I�M ��L�I@M9���   ����   A��=9  ��
H��$�   �������$�   ��$�   �����@ @��E1�L��A������H��$�   �A@ H��$�   Ǆ$�   ����fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$0	   �D$(   �����H��$�   �O�����E1�L��A�щ�������E1�L��A�щ�����H��PH���tH��$�   �_���HǄ$�       1��L���L���{��I�E �+   L���P0�����L��D$|�{��I�E �-   L���P0D�D$|���������UAWAVAUATWVSH��XH��$�   H�EXI�xI�I�YH�M H���   L�uHH�}�M�(�}�H�U�H�U���� I��H�EPH��   H����k���H�U�D�E�H)ă��L�d$ @��M��@��@ ���  ���A��H����D ���  D��@8���  1�1�1�A���A��M��A��E ��(  E��H�}� ��D ���   D��A8���       �   M��t	E���  E��H����   1�E1�� I��H��H9�s1H��H92v�I��LcO��E82tIH��E��H9�D�H��H�
r�I9�tZI�EI;E��   H��I�EH��A������<����     H���f.�     H�E�H�HH9H�\  1�A8��?���H����   H97��   H�E`�H�    ����H#E�I	�H�E L�(L�@H�e�[^_A\A]A^A_]�I�EI9E��  E1������fD  I�EI;E�*  D������f�     I�E L���PP�*���H���w���H97t
H9w�h���Ic$��+UPH��H;MPC�H�U@��Q���@��E����  H�uPH���  1�L�m�1�E��D�}�M��I��L��D�E�� H�H���PD8�tH��H9�tI���D8�u�C�<�H��I��H9�u�L��1�1�L�m�H��M��D�E�D�}������L���$< H��   H�������H)�H��H�D$ H�E�H�ƐIc�I������H��H��H9�u�H�}�A������   �V���H�BH9B�%  1��2���1�I�EI9E�	���I�E H�U�L��L�U�D�E��PHD�E����L�U�H�U��������E1�1������fD  I�E L��D�E�D�U�D�M��PHD�M��    ����    D�U�LD�D�E�DE������H��H� D�E�D�U��U�D�M��PH�U�A�    ����    D�M�HEE�D�U�AE�H�E�D�E�����I�E D�E�L���PHA�����D�E����DEظ    LD�����I�EI;EsPD������1�1��#���H�H��L�U�D�E�H�U��PHH�Uȹ    ����    D�E�E�L�U�HE�H�E������I�E L�U�L��D�E��P�       HA�����L�U����D�E�DEȸ    LD��~���������������AWAVAUATUWVSH���   I�@I�yH��$h  I�H�D$X��M�)H��$P  H��$0  H��$8  H�|$`��$�   H�   H��H��$�   �� H;�$p  I��H��$X  �     �\  L��$p  ���H�e  @��H��$�   f�     ���A��H��A��E ��*  E��M����@ ���  ��D8���  D�>G��<9  L��E��u'I�$L�J@H��w��I9��o  ��tC��<9  A��A��%�6  I�T$0��B ��  H��t	E����   ��I�$D�T$p��L���P �L��A��I�$�P D8�t<H��tD�T$pE����   ��I�$��L���P�L��A��I�$�PD8��5  H�CH;C�s  H��H�CH�������I9�tH��$X  � ���������H�    ����H#l$XH	�H��$0  H�H�hH���   [^_]A\A]A^A_�@ H�CH;C��  �����f.�     H�CH;C��  ��3���f.�     L�~M9��w  D�^G��9  M��E��u,I�$H�Bv��H�@@H9��e  E����  G��9  E��A��E�g  A��O�]  A��E��E1�E1�H��$8  D��$�   D�L$xD�D$pH� H�@@H;�$�   �Q  H�t$X��H�    ����H��$�   H!�H#l$`H	Ƌ�$�   H�t$XH	�H�l$`��� H��$X  D�D$pD�L$xD��$�   �    �x8 �W  D�H^E��D��$�   �!  D��$�   Ƅ$�    H��$�   H��$8  H��$�   H�D$8H��$`  H��$�   L��$�   H��$�       �   L��$�   H��$�   L��$�   H�D$0H��$X  H�D$(H��$P  H�D$ �������$�   H�    ����H��$�   H!�H	փ����H��@��H����@ ��N  M��t@��uV��@8�uH��$X  �H�D$hH��$�   H�    ����H!�H#t$XH	�H�D$hH��$�   ��H	�H�t$X��I�w�,���1�I�MI9Mr�I�E L���PH������H�FI9��  �NH���J u�@ ��B t	H��I9�u�E1�A���VfD  D��M����@ �uq��@8�tH��t	E���}   D��I�T$0���B t`H�CH;C��   H��H�CA�����A���A��H��@��D �t�H�CH9C��  1�M����@ �t�I�EI9E��  1�@8�u�D���2���@ H�CH;C�"  �I�T$0�J ���������I�EI9E��  1�D8�����H��$X  �    �����H�CH9C�?  E1������f�     H�H���PP�,���f�L�~M9���  �vE��A��49  I������  I�$H�|r��@��H�@@H9��>  E���b���E��49  �U���D  D�T$pA��E1�L��A��D�T$p�t��� D��$�   D��$�   Ƅ$�    ����� H��D��$�   D��$�   D�D$xH�D$p�~o��H�D$pD�D$xD��$�   D��$�   H�L�Z0H��q��I9��X���D�T$x�%   H��D�D$pA��D�T$xA��D�D$p�/����E1�1�E1����� H��$�   H��$`  H�    ����H�t$X�T$8L��$�   D��$�   L��$�   D�\$@H��$8  H�\$0H��$X  H!�H#L$`H	�H�t$XH�\$(H��$P�         L	�H��$�   H�L$`L��$�   I��L��$�   H��$�   H�\$ ��H��$�   H��$�   H�D$h���N���H�D�D$xH��D�L$p�PHD�L$p����    D�D$xAE�HD������I�E D��$�   L��T$xD�L$p�PH�T$x����    D�L$pLD�D��$�   AE�����f.�     1�H�HH9H�����H� �T$pH���PH�T$p����    HD�D��|���f.�     H�H��D�D$p�PH�    D�D$p���HD��2�����A��������L�\$xA��E1�L��D�L$p��L�\$xA��D�L$p�r����    H�H���PP����H�D�T$pH���PH�    D�T$p����    DE�HD��^���I�E L��D�T$x�T$p�PH�T$p�    ����    D�T$xLD�E��8���D��$�   E1�L��D�T$xD�L$p��D��$�   ��D�T$xA��D�L$p����L������H��$X  �    �����H�D�T$pH���PH�����D�T$p���Eи    HD��(���H�H���PH��������Eи    HD��C�������������AWAVAUATUWVSH��   H�I�(I�XM�!H�@@I��H��H�  M�qD��$(  ��$0  H9���  H��$  H���   �_� H��$  �    �x8 �  �P^@����$�   �3  D��$�   Ƅ$�    H��$�   L��H�l$pH�D$8H��$   L�L$`H��$�   H�\$xL�D$pL�d$`L�t$hH�D$0H��$  H�D$(H��$  H�D$ ������$�   H�    ����L��$�   H!�H	Ã��@��M����@ �A���I  A�����M��t���  @8�uH��$  �L�>H�^H��H���       �   [^_]A\A]A^A_��    H��H�D$X�j��H�D$XH��l��H�L�J0�%   I9�������%   H��A�щ�����@��$�   D��$�   Ƅ$�    ����� D��E��L�d$pL��H��$   D�D$@L�L$pH��$�   L��$�   H��$�   L�t$xH�|$0H��$  D�|$8H�|$(H��$  H�|$ ������fD  1�I�|$I9|$�����I�$L���PH����������f�     1�I�GI9G�����I�L���PH����    AD�LD�������AWAVAUATUWVSH��   H��$   M�0I�XI�9H��I��I�iH���   D��$  D��$   ��� H��$  �    �x8 �  �P^E�䈔$�   ��   D��$�   D��$�   Ƅ$�    H��$�   L��L�t$`H�D$8H��$  H�L$pL�L$PH�\$hL�D$`H�|$PH�l$XH�D$0H��$  H�D$(H��$   H�D$ �����D$xH�    ����L�t$pH!�H	Ã��A��M����D �A����   �����H��t����   A8�uH��$  �H��L�6H�^H�Ę   [^_]A\A]A^A_�D��$�   Ƅ$�    ����f.�     H��H�D$H��g��H�D$HH�j��H�L�B0�%   I9�������%   H��A�Љ�����E1�I�FI9F�O���I�L���PH����    ED�LD��1����1�H�OH9O�3���H�H���PH���������������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$�       PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[ÐH��  H�H�@H9�u1��f.�     H���������������AVAUATUWVSH��   H��$�   �AoI�)M�qI��H��)L$@L��$�   H���   ��� foT$@H��H�l$`H�@L�L$`L�t$hH��$�   )T$pL�D$pH�@H�\$ L�l$(H�D$8H��$   H�D$0��  H��$�   H�D$@foD$@fĄ$�   )D$P�D$XH�|$Pfo\$Pf���)\$@��H���� ؉�u_fA�����H���t��u.8�uA�M H�|$@fod$@L��A$$H�Đ   [^_]A\A]A^�H�EH;EsD� f�������     H�GH;Gs6� f����    �    D�HD��z���f�     H�E H���PH�@ H�H���PH�����AVAUATUWVSH��   H��$�   �AoI�)M�qI��H��)L$@L��$�   H���   �l� foT$@H��H�l$`H�@L�L$`L�t$hH��$�   )T$pL�D$pH�@ H�\$ L�l$(H�D$8H��$   H�D$0�i  H��$�   H�D$@foD$@fĄ$�   )D$P�D$XH�|$Pfo\$Pf���)\$@��H���� ؉�u_fA�����H���t��u.8�uA�M H�|$@fod$@L��A$$H�Đ   [^_]A\A]A^�H�EH;EsD� f�������     H�GH;Gs6� f����    �    D�HD��z���f�     H�E H���PH�@ H�H���PH�����AVAUATUWVSH��   �AoI��       )M�qL��$  H��$�   I��H�D$8   H�D$HH��$  H��$�   �D$0'  L�L$p�D$(    L��$�   )L$PH�D$@H��$�   H�D$ Ǆ$�       )�$�   H�l$pL�t$x�  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   ��$�   D�Ad�ɍ�����H��$   AHЉQf�����H���� ؉�uqfA�����H���t��u.8�uA�M H�|$Pfod$PL��A$$H�İ   [^_]A\A]A^�H�EH;EsV� f�����8�u��fD  A�M �f�     H�GH;Gs6� f����    �    D�HD��h���f�     H�E H���PH�@ H�H���PH�����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[Ð1�Ð������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[ÐAWAVAUATUWVSH��HA�
   I�@I�qI�M�!H�D$0��H��$�   H��$�   H���   ��� H��$�   I��tH��$�   A��  �   AD�A��f�����L�d$(@��1�E1�H��A��L��A���   H�|$( D����D ���   H;�$�   D���&  @8��  H��t	E���.  A��H�>A�*   H���W`�PЀ�	�@  C����D�|P�D��A��;�$�   �   D�;�$�   �  �����A��H�CA��A��H;C��   H��H�CH��A�����fA���A��H��@���       D ��,���H�CH;C�  � f����    �    HD�E�H�|$( ��D ��	���H�L$(H�AH;A��   � f����    �    E�HEL$(H;�$�   H�L$(�����H��H;�$�   D��uFH��$�   D�8�Yf�H�CH;C��   �f����    HD�����H�H���PP����H��D��H��$�   u?H��u9H��$�   E�W�D�H��$�   f�l$0H�t$0H�H�pH��H[^_]A\A]A^A_�H��$�   ���f�H�D�D$>H���PHD�D$>������    H�L$(D�D$?�T$>H��PHD�D$?�T$>�����H�H���PH���,��������������AVAUATUWVSH��   H��$�  �AoI�)M�iI��H��)L$PL��$�  H���   �<� foT$PǄ$�       H��$�   H�@L�L$pL��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$   H�PxH��$  H���   H���   )�$�   H��$  H��H��$  H��$�   H�l$pH�D$@H��$�   H�D$(H��$�   H�D$ H�\$8H�D$0   L�l$x��  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   H��$�  ��$�   �Jf�����H���� ؉�uufA�����H���t��u28�uA�$H�|$Pfod$PL��A&H��   [^_]A\A]A^�D  H�EH;EsV� f������f.�     A�$�f�     H�GH;G�       s6� f����    �    D�HD��d���f�     H�E H���PH�@ H�H���PH�����UAWAVAUATWVSH��hH��$�   H�EhL�m`�Ao �Ao	H�M0H�]XH���   )E�)M��J� I��J��   H���膹��H�U�H)�H�E�H�U�H�E�L�|$ H���J����t$H�Ep�H�E0foU�H�e�[^_A\A]A^A_]��U�H�M���J��M���t�1�E1�� I�$L���P0f9�tH��I9�tH���f9�u�C�4�H��I��I9�u�1�I���  Ic7A�   H����c��I��f.�     Kc�H����c��I9�LG�I��M9�r�H�M�H�AH;A�  H��H�AH�������L9�f�U�����H�M�A�   H��tH�AH;A�  � E1�f�����  f�}��H�M���H���� �A���m  A8������L�?E1���    I��C��M9�C��v2Kc4�H�M�H��H��B�4�E�t
f�����   f9�u�I��M9�w�I�������I���W���H�M�H�AH;A��  H��H�A�����H��f�E�IcH�4�I��H���b��H9�H���9  A������6fA9�� ���H�M�H�AH;A�
  H��H�AH��fD�e�H9���   H�U�H�M���G���������H�M�D�4~�E�H��t�f���u�H�AH;A��   � f���u�H�E�    �y���D  H�AH;AsF� f��������H�E�    �����H�AH;AsP� 1�f����z���H�E�    D���j��� H�L�M��PHL�M��H��PP�����H�E�    A�   ����H�D�]��PHD�]��H��PH�����H��PP�����H9������H��       EPD�(�����H��PH�#���H��PP�q���AVAUATUWVSH��p  H��$�  �AoI�)M�iI��H��)L$PL��$�  H���   �� H��$�   H�@L�L$pL��$�   H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$�   H��P  H��$�   H��X  H��$�   H��`  H��$�   H��h  H��$�   H��p  H��$�   H��x  H��$   H���  H��$  H���   H��$  H���   H��$  H���   H��$   H���   H��$(  H���   foT$PǄ$�       H��$0  H���   H��$8  H���   H��$@  H��   H��$H  H��  H��$P  H��  H��$X  H��  H��   H�\$8H�D$0   )�$�   H��$`  H��H��$h  H��$�   H�D$@H��$�   H�D$(H��$�   H�D$ H�l$pL�l$x�  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   H��$�  ��$�   �Jf�����H���� ؉�upfA�����H���t��u-8�uA�$H�|$Pfod$PL��A&H��p  [^_]A\A]A^�H�EH;EsV� f������f.�     A�$�f�     H�GH;Gs6� f����    �    D�HD��i���f�     H�E H���PH�@ H�H���PH�����AWAVAUATUWVSH��H  L�5; E1�H��$�  H��$�  �Ao�AoH���   H��$�  H��H��$�  )�$�   )�$�   �J� H��H�D$X��� H��H���j]����$�   Ǆ�       $�       H��$�   I��H��$�   H�D$`f���@��H����@ ����n  f��$�   �H��$�   ��H���� Љ���   @8׋�$�   ��   M9���   ����   H�K�,$E1�H��L�,.A�U I�|$�P`<%uGH�E1�H���T.�P`Ǆ$�       <E�  <O�  ��A<8�I  ��Ic�L���@ H��$�   A�m ��$�   H��t
f����=  f9��c  ��$�   I����$�   �����H�AH;A�   � 1�f��������ꋄ$�   HǄ$�       @8�����M9�u��tH��$�  �H��$�  fo�$�    H��H  [^_]A\A]A^A_�@ H�AH;A��  � 1�f����u���HǄ$�       ���b���H�I�|$E1�H���T.�P`�����D  ��$�   H�L$`��A��E1�H����H��P`<	�"  ��$�   ��$�   �    L�gH��$�   �����H�AH;A��  � f�����  f9�H��$�   ����� H�AH;A�n  H��H�A�����I�������f��$�   �y���H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@H�D$8@ H��$�  L��$�   H��$�  L��$�   H�D$0H��$�   H�D$(H��$�  H�D$ �L���H��$�   ��$�   H��$�   f��$�   ������    H�D$XH��$�   fo�$�   fo�$�   H�@H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$   H���   H��$  H���   )�$�   )�$�   H��$  H��$�   H��$�  H�D�       $0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ����H��$�   ��$�   H��$�   ��$�   f��$�   ���������$�   H��$�  �A���� H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   H��$  H��   H��$  H��  H��$   H��  H��$(  H��  H��$0  H��   )�$�   )�$�   H��$8  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ����H��$�   ��$�   H��$�   ��$�   f��$�   ���@�����$�   H��$�  �A�)���f�     H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0'  L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ������$�   H��$�   ��$�   ��H��$�   f��$�   �j�����$�   D�Ad�ɍ�����H��$�  AH��A�C��� H�L��3 H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   H�l$8����H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(    H��$�  H��$�   H�D$ L��$�   L��$�   �������$�   H��$�   ��$�   ��H��$��          f��$�   �7�����$�   H��$�  �A� ���H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(   �.���H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0;   L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ����D��$�   H��$�   ��$�   E��H��$�   f��$�   ������$�   H��$�  �A�����H�L�B1 H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   �����H��$�   H��$�  H�D$8   H�D$HH��$�  L��$�   H��$�   �D$0<   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ����D��$�   H��$�   ��$�   E��H��$�   f��$�   �������$�   H��$�  ������f�H�L�,0 H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   ����f�H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@ H�D$8�������$�   H�L$`��8��L��   H��D��A�Q�������H��$�  L��$�   H�D$0   H��$�  H��$�   M��fo�$�   L��$�   H�l$@fo�$�   H��$�   L�l$ H�D$8H��o L��$�   H�L$p)�$�   )�$�   H�D$(L�D$h����H��$�   H��$�   H�L$`H��$�   ��$�   f��$�   � 7���       ��$�   ���@�����$�   �$�   �,���H�L$`��7���-   H��f�D$~H��PPf9D$~t0��$�   H�L$`�7���+   H��f�D$~H��PPf9D$~�����H��$�  M��H�l$Hfo�$�   �D$0   L�D$hL�l$ H��$�  )�$�   H�L$pH�D$@fo�$�   �D$(    H�D$8   )�$�   �����H��$�   H�l$HM��H��$�  L�l$ L�D$hH�D$8   H�L$p�D$0;   H��$�   ��$�   fo�$�   �D$(    )�$�   f��$�   H��$�  fo�$�   )�$�   H�D$@�`���H��$�   ��$�   H��$�   f��$�   ����H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   )�$�   )�$�   H��$  �����f.�     H�D$XH��$�   fo�$�   fo�$�   H�@H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$   H��P  H��$  H��X  H��$  H��`  H��$  H��h  H��$   H��p  H��$(  H��x  H��$0  H���  )�$�   )�$�   H��$8  �[���@ H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@0H�D$8����H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ������       H��$�   ��$�   H��$�   ��$�   f��$�   ���)�����$�   H��$�  �A����f���$�   H�L$`�3��L��    H��D��A�Q���  H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(
   H��$�  H��$�   H�D$ L��$�   L��$�   �����H��$�   D��$�   H��$�   ��$�   E��f��$�   ��$�   �#����������$�   H�L$`��2��E1�H����H��P`<
�����H��$�   �8 A����������fD��$�   �����H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �����D��$�   H��$�   ��$�   E��H��$�   f��$�   ������$�   H��$�  ���A�����H��PH�����f�H��PH�f���D  HǄ$�       1�����H��$�   A������
 H��$�   fD��$�   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$0	   �D$(   �����H��PH�f���H��PPH��$�   �����UAWAVAUATWVSH��XH��$�   H�EXI�I�pI�YH�M H���   L�uHM� H�U�H�u�f�u�H�U�蒭 I��H�EPH��   H����ʞ��H�U�H)�f���L�l$ @��M��@��@ ��J  f���A��H����D ��  D��@8���  1�1�1�f�}��A��M��A��E ��D  E��H�       �}� ��D ���   D��A8���   M��t	E���F  �E�H����   L�61�E1��I��H��H9�s4H��H91v�M�D� McO��fC9tHH��E�T� H9�E�L��L�r�I9�tpI�D$I;D$��   H��I�D$�����H��f�E��0���H����    H�M�H�AH;A�~  � f����    �    E�HEM�A8�H�M��$���H����   H97��   D  H�E`��E�f�E�H�E H�u�L� H�pH�e�[^_A\A]A^A_]ÐI�D$I;D$��  � f����    �    LD�DE�����f�I�D$I;D$��  � f����    LD�����I�$L���PP�����H���b���H97t
H9w�S���IcM ��+UPH��H;MPC�H�U@��<����E�@������  H�uPH���  1�L�e�1�M��D�}�M��I��H����I�$L���P0f9�tH��H9�tI���f9�u�C�|� H��I��H9�u�L��1�1�L�e�H��M��D�}��~���I�D$I;D$��  H��I�D$H��   H����ћ��1�H��H)�H�D$ H�E�H��IcD� I����F��H��H��H9�u�����H�}Ⱦ   f�U�����H�BH;B��   � f����    �    HE�E�H�M������I�D$I;D$��   � 1�f����������E1�1�����I�$D�E�L��D�M��PHD�E�D�M�����H�M�D�E�D�M��U�H��PHD�E�D�M��U��]���I�$L���PH�����I�D$I;D$s]� ��f����    LD��@���1�1��0���I�$H�U�L��L�M��PHH�U�L�M��E���H�L�M�H��H�U��PHL�M�H�U������I�$L�M��       L���PHL�M����I�$L���PP�i��������������AWAVAUATUWVSH���   I�A�Ao(H��$x  M�!H�D$pH��$`  H��$@  )l$PL�l$PH��$H  �l$XH�   H��H��$�   臨 H;�$�  H��H��$h  �     �  H��	  M��H�D$x�   @ H��    H��D��P���  M��t	E���M  ��H�H���P@�H�ى�H��P@f9�t1M��t	E���=  ��H�H���P0�H�ى�H��P0f9��v  I�FI;F�+  H��I�FH�������H9�$�  �]  H��$h  ����K  f���A��M����D ��  D��f�|$p�@��M��A��A ���  A��D8���  H�E1�H����P`<%�����H�~H9�$�  ��  H�E1�H���V�P`D��A��E��  1�E1�A��O��  H��$H  L�t$Pf�l$XH� H�@@H;D$x�/  H�D$pL��$�   H��$�   foT$PH��$�   )�$�   详 H��$h  �%   L� �    H��A�PPE��f��$�   ��  fD��$�   1�f��$�   H��$�   H��$H  H�D$8H��$p  H��$�   fo�$�   L��$�   fo�$�   L��$�   )�$�   H�D$0H��$h  )�$�   H�D$(H��$`  H�D$ ����H��$�   H��$�   H��$�   H��$�   ��$�   f��$�   �'����tH��$h  �H��$�   H��$�   H�wH9�$�  H�D$PH��$�   foD$PfĄ$�   )D$`foL$`H��$�   L�t$`)L$P�l$h�����M��H��$@  L�l$Pf�l$Xfol$P(H���   [^_]A\A]A�       ^A_�H��H9�$�  L��$�  u�#@ H��I9�tH��    H��D��P��u�H��$x  E1���E1�H�݉��jf.�     M��D���� ���   ��@8���   M��t	E����   D��H�E �    H���P����   I�FI;F�-  H��I�F�����f���A��M��@��D �t�I�FI;F�  � f���MD�AE�M���� ��r���I�D$I;D$�  � f���AE�MD�@8��U���f�     H���H��$x  �%���I�FI;F�   D� fA���MD��,���I�D$I;D$�4  � f����    �    DE�LD�D8��3���H��$h  M���    �+���fD  I�FI;F��  � f����    �    LD�E������D  I�L���PP�����f�H�~H9�$�  ��  H�E1�H��fE���V�P`A��D�������fD��$�   1�fD��$�   f��$�   �m���I�FI;F��  �f����    LD������     H�t$pH��$�   �T$@fol$PL��$�   L��$�   D�l$8L��$�   H��$H  )�$�   H��$�   H��$p  H�t$0H��$h  H�t$(H��$`  H�t$ ��H��$�   H��$�   ����fD  I�D�D$`L���PHD�D$`������    I�$D��$�   L��T$`�PH�T$`D��$�   ������    I�L���PHD�������I�FI;Fsy�f����    LD�����I�L���PP�����I��T$`L���PH�T$`����I�$�T$`L���PH�T$`����H��$h  M���    ����I�L���PH���q���I�L���PH���y������       ��������AWAVAUATUWVSH���   )�$�   H��Ao8I�)M�iH�@@I��I��H�e  L��$0  H��$8  ��$H  H9Ћ�$P  �n  I���   )|$Pf��詠 �    �%   L� H��A�PP@��f��$�   �  f@��1�f��$�   f��$�   f��$�   H��$�   L�t$ L��H�D$8H��$@  H��$�   H�t$(L�L$pL��$�   )�$�   H�l$pH�D$0L�l$x����H��$�   H�D$PfoD$PfĄ$�   )D$`�D$hL�t$`foL$`f���)L$P��M���� ؉���   fA�����H���t����   8�u�L�t$PfoT$PA$(�$�   L��H���   [^_]A\A]A^A_�fD  1�f��$�   f��$�   �����f�     @����H�t$(L���|$@H��$@  L��$�   )�$�   L��$�   H��$�   L��$�   �\$8H�|$0L�t$ ���c����     I�FI;FsF� f����    �    D�LD�����f�     H�EH;Es&� f�����������    I�L���PH�D  H�E H���PH�ѐ���AWAVAUATUWVSH��   H��$  �AoI�)M�iI��I��)L$@H��$  H���   ��$(  D��$0  �+� �%   L� �    H��f��A�PPE��f��$�   �  1�f��$�   f��$�   H��$�   foT$@H�t$ L��H�D$8H��$   L�L$`H��$�   H�|$(L�D$p)T$pH�l$`H�D$0L�l$h�,���H��$�   H�D$@foD$@fĄ$�   )D$P�D$XL�t$Pfo\$Pf���)\$@��M���� ؉���   fA�����H���t��u.8�u�L�t$�       @fod$@L��A$$H�Ĩ   [^_]A\A]A^A_�H�EH;Esc� f�������    fE��1�f��$�   fD��$�   f��$�   �����I�FI;Fs1� f����    �    D�LD��V���@ H�E H���PH�@ I�L���PH�ǐ����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[ÐAWAVAUATUWVSH���   H��$`  �Ao �Ao	H���   H��$@  H��)�$�   )�$�   贚 H��� H�D$`�s4��H��H��$`  H���   H�@H��H�3H���]  H�~@ H�FdH�D$P��  �D$ �~  H��$�   HǄ$�       H�D$HH��$�   Ƅ$�    H��$�   tH�L$H�    �ή H��$�   �    HǄ$�       H�AH�L$@H��$�   Ƅ$�    藮 H�Fe1�E1��D$~ H�D$8�F`1��D$x    H�D$X    ��$�   H��$�   H�D$hH�D$h�<(��  �(H�=� Hc�H����    A�   H���P  H�|$X��D!�����  �|$~ ��  L�v8��$�   A�   A�����H��$�   f����@��H��@��@ ���  ��$�   �H��$�   ��H��t���]  1�L;d$X��	  @����	  H��$�   ��$�       �   H��t	�����  C8&��  H��$�   H�AH;A�I	  H��H�AD��$�   I��D���Z���f.�     ��$�   A�����H��$�   �   fD  H��Q H+D$PH��$�   H�L�gD�,H�T$@H��$�   H��H9���  H��$�   I9��u  D�,8H��$�   ��L��$�   �D8 H��$�   H�AH;A��  H��H�AǄ$�   ������������@��H��A��A ���  ��$�   �H��$�   ��H��A��A ��c  @8��H	  ��$�   H��$�   ���u	H����  H�L$8@��A�
   �5��H�������@8~!A��E��   �F ���>  @8~"�1  E���:  ���:  H�T$HH��$�   H��$�   H��H9�L�g��  H��$�   I9��o  �8H��$�   1�L��$�   �D8 �����H�~@ ��  H�~P L��$�   L��$�   �*  �|$A��A���o  f�     H��$`  �@uRH�|$X@�ǅ���@�u>���
  ��A�   �,  ��$�   <t<�-  �|$ �"  �    H�F0E1�A�����H��$�   H�D$p��$�   ���@��H��A��A ���  ��$�   �H��$�   ��H��t���  1�L;l$p��@ ���  ��$�   H��$�   ���u	H����  H�V(B8*��  H��$�   H�AH;A��  H��H�AD��$�   I��D���Y����     L��$�   L��$�   L��L���E������  E1�H���������$�   A�����H��$�   �   fD  ��$�   �H��$�   ��H��A��A ����         @8���  ��$�   H��$�   ���u	H���h  H�|$`��H�W0�B ��  H��$�   H�AH;A�  H��H�AD��$�   D�����@��H��A��A ��a���1�H�AH9A�Q���H��PH����B���HǄ$�       D���.���1�H�AH9A�����H��PH1҃���|���HǄ$�       D���h���f�     1�H�AH9A�,���H��PH�������HǄ$�       D���	���H�AH;A�?  �8�<����    H�L$@E1�E1�H��H�D$    脫 H��$�   �b����    H�L$HE1�E1�H��H�D$    �T� H��$�   �h����    �   ����fD  H��PPH��$�   �B����FX����  �\$xA�   1�������   ����A��H��$�    ��   H��$h  �H��$�   H��$�   ������tH��$h  �H��$@  fo�$�   H��$�   H�D$@H��H9�t�� H�D$HH��$�   H��H9�t�� H��$@  H���   [^_]A\A]A^A_�H�AH;A�  H�|$`D� H�W0B�B �����f�     D����E�������@�������H�D$hH���<(�W���1�A�   ���     1�H�AH9A�����H��PH1҃�������HǄ$�       D�������H�~P �D$�8���H�AH9A�����H��PH�����1׃�������HǄ$�       �o���fD  L�vH�
����    ��$�   L�����H�T$`��H�R0�B �����H��$�   �.� Ǆ$�   ����A�   �����     L��$�   L��$�   L��L�����       �������   H�~P udH�~@ �/���1�A�   �D$~�����    H�AH9A�����H��PH�����1׃�������HǄ$�       ����f.�     L��L���u��������  H�~@ �����H�~P ������w���1�H�AH9A����H��PH�������HǄ$�       �������H�AH;A��  �8C8<&�M����
���1�H�AH9A�����H��PH��������HǄ$�       D�������H�AH;A��  H�V(B�*8�(���M�������H��$`  �@�D$p%   A��@���X���f�H��PPH��$�   �����H��PPH��$�   ����f.�     L;d$X�Q���H��$�   �&  �|$~ t*H��$�   �80tH�L$@A�   E1�1��D$ -   蕐 H��$�    t:�D$x��E��H�|$HE�H���?� H�VI��H�N�Oi ��uH��$h  �E��t	9^X�����H�T$@H��$p  �Б ����H��PPH��$�   �����     H��PH����������HǄ$�       D�������E1��     H��$�    A�   �G�������fD  L;l$p�y���A�   �����f.�     H�L$@E1��0   �>V��H�������H���L��$�   �  H�L$@L9�LF�1�耣 ������$�   L���l��H�V88�����H�F@H��$�   H�D$X�� Ǆ$�   ����A�   �Z�����$�   L���%��H�VH8�����H�FPH��$�   H�D$X�S� A�   �D$~Ǆ$�   ���������     �p   膻 H���@    1�H��N f�V H��H��H�F    H�       �F    H���F" H�H�F(    H�F0    H�F8    H�F@    H�FH    H�FP    H�FX    �F`    �Fo ��' H��$`  H��I��H���   �Z H�3�����@ E�������H��$�   �2����S����|$@���%�����$�   ������$�   �9�������H��PH����^���HǄ$�       �M���H��PH����/���HǄ$�       ����E�������E1������H��PH����-���HǄ$�       ����I�@�H���tH���{��������H��$�   �  �f���H����� H�H���P�� H���޻ ��H����� H�������H��H�D$@H��$�   H��H9�t�n� H�D$HH��$�   H��H9�t�S� H��軀��H���ؐ�����AWAVAUATUWVSH���   H��$`  �Ao �Ao	H���   H��$@  H��)�$�   )�$�   �Ċ H��� H�D$`�$��H��H��$`  H���   H�@H��H�3H���]  H�~@ H�FdH�D$P��  �D$ �~  H��$�   HǄ$�       H�D$HH��$�   Ƅ$�    H��$�   tH�L$H�    �ޞ H��$�   �    HǄ$�       H�AH�L$@H��$�   Ƅ$�    觞 H�Fe1�E1��D$~ H�D$8�F`1��D$x    H�D$X    ��$�   H��$�   H�D$hH�D$h�<(��  �(H�=� Hc�H����    A�   H���P  H�|$X��D!�����  �|$~ ��  L�v8��$�   A�   A�����H��$�   f����@��H��@��@ ���  ��$�   �H��$�   ��H��t���]  1�L;d$X��	  @���       ��	  H��$�   ��$�   H��t	�����  C8&��  H��$�   H�AH;A�I	  H��H�AD��$�   I��D���Z���f.�     ��$�   A�����H��$�   �   fD  H�	B H+D$PH��$�   H�L�gD�,H�T$@H��$�   H��H9���  H��$�   I9��u  D�,8H��$�   ��L��$�   �D8 H��$�   H�AH;A��  H��H�AǄ$�   ������������@��H��A��A ���  ��$�   �H��$�   ��H��A��A ��c  @8��H	  ��$�   H��$�   ���u	H����  H�L$8@��A�
   �%��H�������@8~!A��E��   �F ���>  @8~"�1  E���:  ���:  H�T$HH��$�   H��$�   H��H9�L�g��  H��$�   I9��o  �8H��$�   1�L��$�   �D8 �����H�~@ ��  H�~P L��$�   L��$�   �*  �|$A��A���o  f�     H��$`  �@uRH�|$X@�ǅ���@�u>���
  ��A�   �,  ��$�   <t<�-  �|$ �"  �    H�F0E1�A�����H��$�   H�D$p��$�   ���@��H��A��A ���  ��$�   �H��$�   ��H��t���  1�L;l$p��@ ���  ��$�   H��$�   ���u	H����  H�V(B8*��  H��$�   H�AH;A��  H��H�AD��$�   I��D���Y����     L��$�   L��$�   L��L���U������  E1�H���������$�   A�����H��$�   �   fD  ��$�   �H��$�   �       ��H��A��A ���  @8���  ��$�   H��$�   ���u	H���h  H�|$`��H�W0�B ��  H��$�   H�AH;A�  H��H�AD��$�   D�����@��H��A��A ��a���1�H�AH9A�Q���H��PH����B���HǄ$�       D���.���1�H�AH9A�����H��PH1҃���|���HǄ$�       D���h���f�     1�H�AH9A�,���H��PH�������HǄ$�       D���	���H�AH;A�?  �8�<����    H�L$@E1�E1�H��H�D$    蔛 H��$�   �b����    H�L$HE1�E1�H��H�D$    �d� H��$�   �h����    �   ����fD  H��PPH��$�   �B����FX����  �\$xA�   1�������   ����A��H��$�    ��   H��$h  �H��$�   H��$�   ������tH��$h  �H��$@  fo�$�   H��$�   H�D$@H��H9�t�ư H�D$HH��$�   H��H9�t諰 H��$@  H���   [^_]A\A]A^A_�H�AH;A�  H�|$`D� H�W0B�B �����f�     D����E�������@�������H�D$hH���<(�W���1�A�   ���     1�H�AH9A�����H��PH1҃�������HǄ$�       D�������H�~P �D$�8���H�AH9A�����H��PH�����1׃�������HǄ$�       �o���fD  L�vH�
����    ��$�   L�����H�T$`��H�R0�B �����H��$�   �>� Ǆ$�   ����A�   �����     L��$�   �       L��$�   L��L����������   H�~P udH�~@ �/���1�A�   �D$~�����    H�AH9A�����H��PH�����1׃�������HǄ$�       ����f.�     L��L�����������  H�~@ �����H�~P ������w���1�H�AH9A����H��PH�������HǄ$�       �������H�AH;A��  �8C8<&�M����
���1�H�AH9A�����H��PH��������HǄ$�       D�������H�AH;A��  H�V(B�*8�(���M�������H��$`  �@�D$p%   A��@���X���f�H��PPH��$�   �����H��PPH��$�   ����f.�     L;d$X�Q���H��$�   �&  �|$~ t*H��$�   �80tH�L$@A�   E1�1��D$ -   襀 H��$�    t:�D$x��E��H�|$HE�H���O� H�VI��H�N�_Y ��uH��$h  �E��t	9^X�����H�T$@H��$p  ��� ����H��PPH��$�   �����     H��PH����������HǄ$�       D�������E1��     H��$�    A�   �G�������fD  L;l$p�y���A�   �����f.�     H�L$@E1��0   �NF��H�������H���L��$�   �  H�L$@L9�LF�1�萓 ������$�   L���|���H�V88�����H�F@H��$�   H�D$X�� Ǆ$�   ����A�   �Z�����$�   L���5���H�VH8�����H�FPH��$�   H�D$X�c� A�   �D$~Ǆ$�   ���������     �p   薫 H���@    1�H��> f�V�        H��H��H�F    H�F    H���F" H�H�F(    H�F0    H�F8    H�F@    H�FH    H�FP    H�FX    �F`    �Fo �� H��$`  H��I��H���   �J H�3�����@ E�������H��$�   �2����S����|$@���%�����$�   ������$�   �9�������H��PH����^���HǄ$�       �M���H��PH����/���HǄ$�       ����E�������E1������H��PH����-���HǄ$�       ����I�@�H���tH���{��������H��$�   �  �f���H���� H�H���P覲 H���� ��H���� H���q��H��H�D$@H��$�   H��H9�t�~� H�D$HH��$�   H��H9�t�c� H����p��H���ؐ�����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����AWAVAUATUWVSH��   )�$�   H��$  I�8M�h�Ao9H��I��D��$  H���   ��y H�\$pH�|$PL��Ƅ$�    H�L$`I��H�CE��L�l$XH�D$pH��$   L�L$@H�D$x    L�D$P)|$@H�\$0H�D$(H�t$ tx����H�    ����H�D$`H�T$hL!�L�l$xH��H�D$`H�T$h�D$hH	�M��uNH�L$pH��H�} H�uH9�t�s� �(�$�   H��H�Ĩ   [^_]A\A]A^A_� �����f�       �     H��$(  E1�L���=� H��$(  L�t$pL�8A�D$8<t��t/I�$H�D��H�@8H9�u+M��L��L���]���Z����     L����
����fD  M��L��L��O�.���.���H�L$pH��H��H9�t覦 H���n����������������AUATUWVSH��   I�0M�hM�QH��$  M�	H��HǄ$�       L��$  H��$�   Ƅ$�    ��$    H�KH�t$PH��$�   L�L$@H�L$`L�l$XL�L$@L�T$HL�D$PH�\$0L�d$(H�D$ ��   ����H�    ����H�D$`H�T$hL!�H��H�D$`H�T$h�D$hH	��_ H��$�   L�L$xM��H�D$xH��$  H���=F H��$�   H�u H�}H9�t胥 H��H�Ĩ   [^_]A\A]��;����s���H��$�   H��H��H9�t�M� H���l�������AWAVAUATUWVSH���   H��$`  �Ao �Ao	H���   H��$@  H��)�$�   )�$�   �$w H�� H�D$`���H��H��$`  H���   H�@H��H�;H����  H�@ H�GdH�D$P�	  �D$ �  H��$�   HǄ$�       H�D$HH��$�   Ƅ$�    H��$�   tH�L$H�    �ފ H��$�   �    HǄ$�       H�AH�L$@H��$�   Ƅ$�    觊 H�GfE1�E1��D$~ H�D$8�G`1��D$x    H�D$X    ��$�   H��$�   H�D$hH�D$hB�< ��  B� H��� Hc�H���   I���2  H�|$X��!����  �|$~ �  L�8��$�   A�   A�����H��$�   �   f�f��$�   �H��$�   ��H��@��@ ���       �  8���  L;d$X��  H��$�   ��$�   H��t
f����S	  fC9g�H  H��$�   H�AH;A�
  H��H�AfD��$�   I��D��f�����H��@��@ ��Z���H�AH;A�!  � 1�f����=���HǄ$�       ���*�����$�   H�_zH��$�   fD  f���@��H��A��A ��8  f��$�   �H��$�   ��H��A��A ��4  @8��`  H��$�   ��$�   H��t
f����  H�T$8�    f9��  H��H9�u�f9G"��D���  �o @���n  f9G$�  E���b  ���L  H�L$HH��$�   H��$�   H�QH9�L�u�o  H��$�   I9���  @�4(H��$�   1�L��$�   �D( H��$�   H�AH;A��  H��H�A����������f��$�   ����H�@ ��  H�P H��$�   L��$�   �7  �\$�݃���  H��$`  �@uKH�|$X��E�����u8A����	  A���   ��  ��$�   <t<��  �|$ ��  H�G01�A�����H��$�   H�D$p��$�   �   f��$�   �H��$�   ��H��A��A ���  H;l$p��1� ���  ��$�   H��$�   f���u	H���  H�W(f9j��  H��$�   H�AH;A�;  H��H�AfD��$�   H��D��f�����H��A��A ��X���H�AH;A�|	  � 1�f����;���HǄ$�       D���'���H��$�   L��$�   H��L����������_  1�I���������$�   A�����H��$�   �   �     f��$�   �       �H��$�   ��H��A��A ��M  8��  H��$�   D��$�   H��tfA����U  H�L$`�    H��P����  H��$�   H�AH;A��  H��H�AfD��$�   D��f�����H��A��A ��Z���H�AH;A��  � 1�f����=���HǄ$�       D���)���f�     H��) H+T$PH�L$@H��$�   H� H��L�uD�<H�QH��$�   H9���  H��$�   I9��b  D�<(H��$�   ��L��$�   �D( �����H�AH;A�I  � 1�f��������HǄ$�       D��@8�������   H��$�    ��  H��$h  �H��$�   H��$�   �������tH��$h  �H��$@  fo�$�   H��$�   H�D$@H��H9�t�i� H�D$HH��$�   H��H9�t�N� H��$@  H���   [^_]A\A]A^A_�f�H�AH;A�^  � 1�f��������HǄ$�       D������H�AH;A�C  � f��������HǄ$�       ���� H�L$@E1�E1�H��H�D$    脆 H��$�   �u����    H�L$HE1�E1�H��H�D$    �T� H��$�   ������    �   �+���fD  H��PPH��$�   ������OX���'  �t$xA�   1������   �������A�D$���_������W���H�D$hI��B�< ����1۽   ��H�AH;A�!  � 1�f��������HǄ$�       D������H�AH;A�  D� fA��������HǄ$�       �}���H�P �D$�����L�H�����H��$�   L��$�   H��L����       ��������F  H�P ujH�@ �(���1۽   �D$~������$�   L���`���H�L$`D���    L�	A�Q�����r���H��$�   ��� �����f��$�   �#���H��L�����������o  H�@ �����H�P ������q���f�H�AH;A�  � 1�f����G���HǄ$�       ��8��9���L;d$X�����H��$�   ��  �|$~ t*H��$�   �80tH�L$@A�   E1�1��D$ -   �m H��$�    t;�D$x@��E��H�\$HE�H���K� H�WI��H�O�[F ��uH��$h  �E��t	9wX����H�T$@H��$p  ��n ����H�AH;A�)  � f��������HǄ$�       ����H�AH;A�?  � 1�f�������H;l$pD��HǄ$�       ��1� �����H;l$p�\���H�������H��$`  �@�D$p%   @��������H�AH;A��  � f��������HǄ$�       �����H��PPH��$�   ����H��PPH��$�   �����H��PPH��$�   ����H��PH����H��PH����H��PH����H�L$@E1��0   �2��H���%���H���L��$�   �3  H�L$@L9�LF�1��� �������$�   L������H�WHf9�t���H�GPH��$�   H�D$X��� A������   �D$~fD��$�   �������$�   L���=���H�W8f9�����H�G@H��$�   H�D$X�� A������   fD��$�   �������   ��� H���@    H��H�+ H�G    H��H�G    �G  H���G"    H�H�G(    H�G0    H�G8 �          H�G@    H�GH    H�GP    H�GX    �G`    �Gz �� H��$`  H��I��H���   �7 H�;�V���@���C���H��$�   ������S����\$���8�����$�   �*�����$�   ����������     H��PH�����H��PH����H��PHD�������H��PH�����H��PH�����H��PH�����1�����������D������H��PH�A���H��PH�|���H��PH����I�@�H���tH�����������H��$�   �  ����E1��8���H��H�D$HH��$�   H��H9�t��� H���]]��H���%� H�H���P�Ǟ H���� ��H��H�D$@H��$�   H��H9�t�试 �H���� H���]���������������AWAVAUATUWVSH���   H��$`  �Ao �Ao	H���   H��$@  H��)�$�   )�$�   �tg H�m� H�D$`�� ��H��H��$`  H���   H�@H��H�;H����  H�@ H�GdH�D$P�	  �D$ �  H��$�   HǄ$�       H�D$HH��$�   Ƅ$�    H��$�   tH�L$H�    �.{ H��$�   �    HǄ$�       H�AH�L$@H��$�   Ƅ$�    ��z H�GfE1�E1��D$~ H�D$8�G`1��D$x    H�D$X    ��$�   H��$�   H�D$hH�D$hB�< ��  B� H��� Hc�H���   I���2  H�|$X��!����  �|$~ �  L�8��$�   A�   A�����H��$�   �   f�f��$�   �H��$�   ��H��@��@ ���  8���  L;d$X��  H��$�   ��$�   H��t
f����       �S	  fC9g�H  H��$�   H�AH;A�
  H��H�AfD��$�   I��D��f�����H��@��@ ��Z���H�AH;A�!  � 1�f����=���HǄ$�       ���*�����$�   H�_zH��$�   fD  f���@��H��A��A ��8  f��$�   �H��$�   ��H��A��A ��4  @8��`  H��$�   ��$�   H��t
f����  H�T$8�    f9��  H��H9�u�f9G"��D���  �o @���n  f9G$�  E���b  ���L  H�L$HH��$�   H��$�   H�QH9�L�u�o  H��$�   I9���  @�4(H��$�   1�L��$�   �D( H��$�   H�AH;A��  H��H�A����������f��$�   ����H�@ ��  H�P H��$�   L��$�   �7  �\$�݃���  H��$`  �@uKH�|$X��E�����u8A����	  A���   ��  ��$�   <t<��  �|$ ��  H�G01�A�����H��$�   H�D$p��$�   �   f��$�   �H��$�   ��H��A��A ���  H;l$p��1� ���  ��$�   H��$�   f���u	H���  H�W(f9j��  H��$�   H�AH;A�;  H��H�AfD��$�   H��D��f�����H��A��A ��X���H�AH;A�|	  � 1�f����;���HǄ$�       D���'���H��$�   L��$�   H��L���������_  1�I���������$�   A�����H��$�   �   �     f��$�   �H��$�   ��H��A��A ��M  8��  H��$�   D���       $�   H��tfA����U  H�L$`�    H��P����  H��$�   H�AH;A��  H��H�AfD��$�   D��f�����H��A��A ��Z���H�AH;A��  � 1�f����=���HǄ$�       D���)���f�     H�9 H+T$PH�L$@H��$�   H� H��L�uD�<H�QH��$�   H9���  H��$�   I9��b  D�<(H��$�   ��L��$�   �D( �����H�AH;A�I  � 1�f��������HǄ$�       D��@8�������   H��$�    ��  H��$h  �H��$�   H��$�   �'�����tH��$h  �H��$@  fo�$�   H��$�   H�D$@H��H9�t蹍 H�D$HH��$�   H��H9�t融 H��$@  H���   [^_]A\A]A^A_�f�H�AH;A�^  � 1�f��������HǄ$�       D������H�AH;A�C  � f��������HǄ$�       ���� H�L$@E1�E1�H��H�D$    ��v H��$�   �u����    H�L$HE1�E1�H��H�D$    �v H��$�   ������    �   �+���fD  H��PPH��$�   ������OX���'  �t$xA�   1������   �������A�D$���_������W���H�D$hI��B�< ����1۽   ��H�AH;A�!  � 1�f��������HǄ$�       D������H�AH;A�  D� fA��������HǄ$�       �}���H�P �D$�����L�H�����H��$�   L��$�   H��L������������F  H�P ujH�@ �(���1۽   �D$~�����       ��$�   L������H�L$`D���    L�	A�Q�����r���H��$�   �� �����f��$�   �#���H��L���W��������o  H�@ �����H�P ������q���f�H�AH;A�  � 1�f����G���HǄ$�       ��8��9���L;d$X�����H��$�   ��  �|$~ t*H��$�   �80tH�L$@A�   E1�1��D$ -   ��] H��$�    t;�D$x@��E��H�\$HE�H���u H�WI��H�O�6 ��uH��$h  �E��t	9wX����H�T$@H��$p  �,_ ����H�AH;A�)  � f��������HǄ$�       ����H�AH;A�?  � 1�f�������H;l$pD��HǄ$�       ��1� �����H;l$p�\���H�������H��$`  �@�D$p%   @��������H�AH;A��  � f��������HǄ$�       �����H��PPH��$�   ����H��PPH��$�   �����H��PPH��$�   ����H��PH����H��PH����H��PH����H�L$@E1��0   �#��H���%���H���L��$�   �3  H�L$@L9�LF�1��Cp �������$�   L�������H�WHf9�t���H�GPH��$�   H�D$X�K� A������   �D$~fD��$�   �������$�   L������H�W8f9�����H�G@H��$�   H�D$X��� A������   fD��$�   �������   �F� H���@    H��H�r H�G    H��H�G    �G  H���G"    H�H�G(    H�G0    H�G8    H�G@    H�GH    H�GP    H�GX    �G`    �Gz ��       	 H��$`  H��I��H���   �k' H�;�V���@���C���H��$�   ������S����\$���8�����$�   �*�����$�   ����������     H��PH�����H��PH����H��PHD�������H��PH�����H��PH�����H��PH�����1�����������D������H��PH�A���H��PH�|���H��PH����I�@�H���tH�����������H��$�   �  ����E1��8���H��H�D$HH��$�   H��H9�t�E� H���M��H���u� H�H���P�� H���_� ��H��H�D$@H��$�   H��H9�t���� �H���U� H���]M���������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����AUATUWVSH���   )�$�   )�$�   H��$(  D��$   �Ao �Ao9H��H��)D$@H���   ��V H��$�   E��HǄ$�       Ƅ$�    H�L$pI��H�CH��$�   ��   H��$0  H�\$0L�L$PH��foL$@H�t$ L�D$`)|$P)L$`H�D$(����H��$�   H�D$pH�T$xH��H�D$@fot$@H�T$xf�t$xH�D$pu{H��$�   H��7H9�t�� �(�$�   H��(�$�   H���   [^_]A\A]�H��$0  H�\$0L�L$PH��foT$@H�t$ L�D$`)|$P)T$`H�D$(�U����R����       H��$8  E1�H���=� H��$8  H��$�   I�$L�	L��L�2�PX�L���H��$�   H��H��H9�t�>� H���J��������WVSH���   )�$�   ��$    �Ao M�QH��$  H��$�   H��)D$@M�	H�KH��$  HǄ$�       H��$�   H�L$pƄ$�    ��   L�L$PL�D$`H�\$0L�L$PH�|$(H�D$ )D$`L�T$X����H�D$pH�T$xH�D$@fot$@H�T$xf�t$xH�D$p�; H��$�   L��$�   I��H��H��$  H��$�   ��" H��$�   6H9�t�&� �(�$�   H��H���   [^_�foT$@L�L$PL�D$`H�\$0L�L$PH�|$(H�D$ )T$`L�T$X�����E���H��$�   H��H��H9�t辁 H���&I��������SH��P�Ao H�H��)D$@E��H��$�   L�D$@H�L$0��$�   �L$(H��$�   H�L$ H���PH��H��P[Ð������������SH��`H��$�   �Ao �(H��)D$PE��H�L$@H�H�L$0��$�   L�D$P�|$@�L$(H��$�   H�L$ H���PH��H��`[Ð�SH��@�D$x�Ao�D$ L�D$0H��E��H��$�   )L$0L�L$pH�L$(H��t�
  H��H��@[��     �+  H��H��@[Ð�UAWAVAUATWVSH��   H��$�   )} ���   �Ao8�E�H���   H�}�I��H���   H��D�M��(H���   �}�H���   �; H����Q H��@I��H�t$0I���S9 �m�A�@   H��H�E �D$     H��H��L�m�L�l$(L��� �}���" ��?~R���E�H�H��H����CC��H)�H�t$0I����8 D�E�L�l$(H��H���m��D$     H�       �E L��� �}��" Hc�E1�H��H�CH��H�E �N A�D$8L�m <t ����   I�$H�����H�@8H9���   I��L��L�������E�)}�L�E�L���}� H�\$(L���   H���   �D$ t8��  H�M H��H9�t��~ H���&; �(} L��H�e8[^_A\A]A^A_]��X   ��fD  L��������\��� M��L��L��M�6���k���H�M H��H��H9�t�~ H���: H����E��H���됐AWAVAUATUWVSH���   I� I�xH��$X  H�D$0��$P  M���   L��H��$0  L��A���D$L�D$n��O H�� H�D$8����I��H���   H�@N�$�I�$H����  L�e �CdH�mA8$�'  �C\��$�   H�C8H�D$XH�C@H�D$@L�L9�v:H�D$8A�$H�H0L���Qu�!f.�     ��QtGH��H9�u�L)�uAH��$0  H�F    D��H�t$0H�xH�0H���   [^_]A\A]A^A_�fD  H��L)�t�L��$�   Ƅ$�    I�EL��L�l$PH�T- H��$�   HǄ$�       �~c �CXA��A)�E����   ��L��$�   DH�H�{ �(  G�6�D$     1�L��Mc��*P L�KIc�L�CL��S"H�D$(H��$�   L�d$ � L��$�   I��L+�$�   M9���  L��$�   �  �CX��L��$�   �7  �FLl$@����   ���L$h��  L��$�   Ƅ$�    I�FL��HǄ$�       K�T- H��$�   �b H�NH��$�   �|$hL�%�� H�L$`��L9���L)�!�H�L$pH�E�T$oH�D$8�} �V  �E Ic�L�����C`H�퉄$�   �$�       ���H�CHI��H�D$XH�CPH�D$@�����f�H�|$@ �  H�D$XL����f ��   �F��   H��������L�C0H+�$�   H�S(I9���   H��� �+ fD  �|$o L��$�   ��  I�EH�D$xH��$�   I�VH9��  H��$�   H9T$x��  �T$nB�(I�EH��$�   H��$�   B�D( �O�    �|$o tA�D$nE1�L��L�L$pH��$�   �D$ ��M �fD  L��$�   H��$�   L���xb H��H9l$8�����H�D$@H��$�   H����   H�L$`H9���   E��H��$�   Hc�uH�L$0I��H��P`H��$�   H9�A��H�\$01�I��D��L9�@��H��$�   A��H��$�   tH����y H�D$PH��$�   H��H9��C����y �9���f�H)��D$LA�    �|$h I�ɉD$ �  1�L����L H�\$`�H���Lk0�9��� H�T$XI��H��������I��H)�H��I9���  L���Ra H��$�   H�L$`H9�������w����    �C!H�L$P�D$`I�EH�D$8H��$�   H�QH9��  H��$�   H9T$8��  �L$`E��H�T$8B�(H��$�   H��$�   � �;  LcCXIc�H��������H+�$�   L�I9���  H�L$P�` L��$�   �$����D$nE1�L��L��L�L$p�D$ ��K �����f.�     �p   �x H���@    L��H�� H�C    H��H�C    �C" H��H�C(    H�1�f�C H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co ��� H���   H��M��� I�$����H�L�       $PIc�M��1�H�D$ �C �CX�%���H��L����J ������CeA��E1�H��$�   Mc�H�L$P�D$ ��J H��������H+�$�   H9���   I��L������H�L$PE1�E1�L��H�D$    ��` H��$�   �(���H�D$    E1�E1�L��L����` H��$�   �����   ������   �����H�(� �S' H�� �G' H�-� H�A� �d- H��� �(' H��$�   I��H��L9�t�v H�T$PH��$�   H��H9�t�dv H����=��H����H���x H�H���P�1 H���yx ��H���z H���=���������AWAVAUATUWVSH���   I� I�xH��$X  H�D$8��$P  M���   L��H��$0  L��A���D$T�D$v�G H�֩ H�D$@�\���I��H���   H�@N�$�I�$H���  L�e �CdH�mA8$�7  �C\��$�   H�C8H�D$`H�C@H�D$HL�L9�v:H�D$@A�$H�H0L���Qu�!f.�     ��QtGH��H9�u�L)�uAH��$0  H�F    D��H�t$8H�xH�0H���   [^_]A\A]A^A_�fD  H��L)�t�L��$�   Ƅ$�    I�EL��L�l$XH�T- H��$�   HǄ$�       �.[ �CXA��A)�E����   ��L��$�   DH�H�{ ��  G�6�D$     1�L��Mc���G L�KIc�L�CL��S"H�D$(H��$�   L�d$ �� L��$�   I��L+�$�   M9��  L��$�   �  �CX��L��$�   ��  �FLl$H����   ���L$p�^  L��$�   Ƅ$�    I�FL��HǄ$�       K�T- H��$�   �5Z H�NH�       ��$�   �|$pL�%m� H�L$h��L9���L)�I��������!�H�L$xH�E�T$wH�D$@�} ��   �E Ic�L����    �C`H�퉄$�   ����H�CHI��H�D$`H�CPH�D$H����f�H�|$H ��   H�D$`L����D^ �   �F�   L�C0L��H+�$�   H�S(I9�v_H�6� �a# ��|$w �T$v�5  �T$ L�L$xE1�L��H��$�   �F �,f��|$w t#�D$v�D$ ��L��$�   H��$�   L���Z H��H9l$@�����H�D$HH��$�   H����   H�L$hH9���   E��H��$�   Hc�uH�L$8I��H��P`H��$�   H9�A��H�\$81�I��D��L9�@��H��$�   A��H��$�   tH����q H�D$XH��$�   H��H9��������q ����H)��D$TA�    �|$p I�ɉD$ ��  1�L���E H�\$h�J���Lk0���� H�T$`I��H��������I��H)�H��I9��1  L���bY H��$�   H�L$hH9�������w����    �C!H�L$X�D$hI�EH�D$@H��$�   H�QH9���  H��$�   H9T$@��  �L$hE��H�T$@B�(H��$�   H��$�   � �&  LcCXIc�H��������H+�$�   L�I9���  H�L$X�X L��$�   ����L����[ �����p   �p H���@    L��H�� H�C    H��H�C    �C" H��H�C(    H�1�f�C H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co ��� H���   H��M���� I�$�<���f�     H�L$XIc�M��1�H�D$ ��; ��       CX����H��L���C �����CeA��E1�H��$�   Mc�H�L$X�D$ ��B H��������H+�$�   H9�w]I��L������H�L$XE1�E1�L��H�D$    �Y H��$�   �A����   �,���H��� � H��� H��� ��% H�c� � H�W� � H��$�   I��H��L9�t��n H�T$XH��$�   H��H9�t�n H���&6��H����H����p H�H���P�w H����p ��H����r H����5���SH��P�Ao H�H��)D$@E��H��$�   L�D$@H�L$0��$�   �L$(H��$�   H�L$ H���PH��H��P[Ð������������SH��`H��$�   �Ao �(H��)D$PE��H�L$@H�H�L$0��$�   L�D$P�|$@�L$(H��$�   H�L$ H���PH��H��`[Ð�SH��@�D$x�Ao�D$ L�D$0H��E��H��$�   )L$0L�L$pH�L$(H��t��
  H��H��@[��     ��  H��H��@[Ð�UAWAVAUATWVSH��   H��$�   )} ���   �Ao8�E�H���   H�}�I��H���   H��D�M��(H���   �}�H���   �o( H���'? H��@I��H�t$0I���#& �m�A�@   H��H�E �D$     H��H��L�m�L�l$(L�}� �}�� ��?~R���E�H�H��H����0��H)�H�t$0I����% D�E�L�l$(H��H���m��D$     H�E L�&� �}��f Hc�E1�H��H�CH��H�E ��c I�M�4L��L��L�M �PX�E�)}�L�E�L���}� H�\$(L���   H���   �D$ t=�8	  H�M H��H9�t��k H���( �(} L��H�e8[^_A\A]A^A_]�D  �       �;   ��H�M H��H��H9�t�k H����' H���3��H���됐�������������AWAVAUATUWVSH���   I� I�xL��$X  H�D$0��$P  M���   L��H��$0  L��@�|$Y�D$\f�D$Z�Z= H�C� H������I��H���   H�@N�,�I�] H����  M�,$�KdI�D$fA9M tx�S\��$�   H�S8H�T$PH�S@H�T$8L�U M�LE M��H��   A�R(L)�I��I��uiH��$0  H�F    @�|$YH�t$0H�xH�0H���   [^_]A\A]A^A_�@ �S`H��H�KP��$�   H�SHH�L$8H�T$PI�ULE��x���@ H��$�   E1�HǄ$�       H�QH�L$HH��$�   H��fD��$�   ��y �CXE��H��$�   A)�E����   ��EH�H�{ �<  H�L$HG�4?I��1�Mc��D$     M���e L�KM�L�C�S$L�t$(H��$�   L�l$ � L��$�   I��L+�$�   I��M9�L���  E1�L��$�   fD��CX���M  �FHl$8��   ���T$`��  L��$�   E1�HǄ$�       fD��$�   I�FL��H�T- H��$�   ��x L�~L��$�   �|$`L�-�� ��I9���!�I�D$�T$gH�D$@L��H)�H�D$hA�<$�t  A�$IcD� L���H�|$8 �Y  H�D$PI�VH��$�   � f�D$pH�EH�D$xH��$�   H9���  H��$�   H9T$x�?  �L$pH�Uf�h1�H��$�   f�Lh��   f.�     �F��   H��������?L�C0H+�$�   H�S(I9���   H�,� � �    �|$g H��$�   �m  H�EH�D$pH��$�   I�V�       H9��?  H��$�   H9T$p��  �L$ZH�Uf�hH��$�   1�f�Th�F�|$g t?�D$ZE1�L��L�L$hH��$�   �D$ �Fc �@ L��$�   H��$�   L����x I��L9d$@�r���H�D$8H��$�   H����   I9���   I�π|$Y Ic�H��$�   uH�L$0I��H��P`H��$�   H9��D$Y1�H�\$0I���D$YL9�H��$�   H��$�   @��tH���f H�D$HH��$�   H��H9�������f ����� M���D$\A�    I)Ƀ|$` �D$ �D  1�L���Fb �K����Hk0�����    H�T$PI��H��������?I��H)�H��I9���  L���w H��$�   I9�������|����C"L�uH�L$Hf�D$@H��$�   H�QH9��U  H��$�   I9���  �L$@E1�E��f�hL��$�   fD�Lh�A  LcCXMc�H��������?K�T} L)�I9��B  H�L$H�w H��$�   �����     �D$ZE1�H��L��L�L$h�D$ �4a ������   �e H���@    L��H��� H�C    H��H�C    �C  H���C"    H�H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz �� H���   H��M��� I�] ����f�     H�L$HIc�M��I��H�D$ 1���X �CXH��$�   ����fD  �CfA��E1�L��H�L$HMcωD$ �2` H��������?H+�$�   I9���   M��L������H��L���` ����H�D$    E1�E1�H��L���Rw H��$�   ����D  H�L$HE1�E1�H��H�D$    �$w H��$�       �   ������    H�D$    E1�E1�H��L����v H��$�   �����f�     �   ����fD  �   �����   ����H��� H�Ʈ � H��� �� H�v� �� H�j� �� H��H�T$HH��$�   H��H9�t�c H���*��H��$�   I��H��L9�t���b ��H���,e H�H���P��k H���e ��H���,g H���4*������AWAVAUATUWVSH���   I� I�xL��$X  H�D$0��$P  M���   L��H��$0  L��@�|$Y�D$\f�D$Z�4 H��� H�������I��H���   H�@N�,�I�] H����  M�,$�KdI�D$fA9M tx�S\��$�   H�S8H�T$PH�S@H�T$8L�U M�LE M��H��   A�R(L)�I��I��uiH��$0  H�F    @�|$YH�t$0H�xH�0H���   [^_]A\A]A^A_�@ �S`H��H�KP��$�   H�SHH�L$8H�T$PI�ULE��x���@ H��$�   E1�HǄ$�       H�QH�L$HH��$�   H��fD��$�   �'q �CXE��H��$�   A)�E����   ��EH�H�{ �<  H�L$HG�4?I��1�Mc��D$     M����\ L�KM�L�C�S$L�t$(H��$�   L�l$ ��� L��$�   I��L+�$�   I��M9�L���  E1�L��$�   fD��CX���M  �FHl$8��   ���T$`��  L��$�   E1�HǄ$�       fD��$�   I�FL��H�T- H��$�   �#p L�~L��$�   �|$`L�-˫ ��I9���!�I�D$�T$gH�D$@L��H)�H�D$hA�<$�t  A�$IcD� L���H�|$8 �Y  H�D$PI�V�       H��$�   � f�D$pH�EH�D$xH��$�   H9���  H��$�   H9T$x�?  �L$pH�Uf�h1�H��$�   f�Lh��   f.�     �F��   H��������?L�C0H+�$�   H�S(I9���   H�l� �� �    �|$g H��$�   �m  H�EH�D$pH��$�   I�VH9��?  H��$�   H9T$p��  �L$ZH�Uf�hH��$�   1�f�Th�F�|$g t?�D$ZE1�L��L�L$hH��$�   �D$ �Z �@ L��$�   H��$�   L���p I��L9d$@�r���H�D$8H��$�   H����   I9���   I�π|$Y Ic�H��$�   uH�L$0I��H��P`H��$�   H9��D$Y1�H�\$0I���D$YL9�H��$�   H��$�   @��tH����] H�D$HH��$�   H��H9��������] ����� M���D$\A�    I)Ƀ|$` �D$ �D  1�L���Y �K����Hk0�����    H�T$PI��H��������?I��H)�H��I9���  L����n H��$�   I9�������|����C"L�uH�L$Hf�D$@H��$�   H�QH9��U  H��$�   I9���  �L$@E1�E��f�hL��$�   fD�Lh�A  LcCXMc�H��������?K�T} L)�I9��B  H�L$H�En H��$�   �����     �D$ZE1�H��L��L�L$h�D$ �tX ������   ��\ H���@    L��H��� H�C    H��H�C    �C  H���C"    H�H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz �� H���   H��M����� I�] ����f�     �       H�L$HIc�M��I��H�D$ 1��6P �CXH��$�   ����fD  �CfA��E1�L��H�L$HMcωD$ �rW H��������?H+�$�   I9���   M��L������H��L���AW ����H�D$    E1�E1�H��L���n H��$�   ����D  H�L$HE1�E1�H��H�D$    �dn H��$�   ������    H�D$    E1�E1�H��L���6n H��$�   �����f�     �   ����fD  �   �����   ����H�� H�� �Y H�¥ � H��� � H��� � H��H�T$HH��$�   H��H9�t�WZ H���!��H��$�   I��H��L9�t��6Z ��H���l\ H�H���P�c H���V\ ��H���l^ H���t!������H��HH�D$xH�D$0H��$�   H�T$0L�D$ H�L$ A��� L�L$(E1�H�D$8� H�T$pH�L$ H�
H��$�   H�L$0H�
H��HÐSH��0H�L$hH�D$pM9�M��M��H�L$ H�D$(t|A����� wuH�\$ �f.�     I��M9�t7A����� w<H���� ��u�H�L$ �   H�T$`L�H�T$xH�
H��0[�H�L$ 1����    H�L$ �   ��@ 1��Ƹ   뿐����WVSH��0H�D$pL�D$ H�X�H��L��L�L$(t?H�|$ f�     ��� H���� =�� ��H����H����u݋D$ )�H��0[^_�1�H��0[^_Ð����H�D$(L� �   Ð�1�Ð�������������   Ð���������1�Ð������������H��XH��$�   H�D$@H��$�   H�T$@L�D$0H�L$0A��� L�L$8A�   �D$     H�D$H�% H��$�   H�L$0�       H�
H��$�   H�L$@H�
H��X�H��HH�D$xH�D$0H��$�   H�T$0L�D$ H�L$ A��� L�L$(E1�H�D$8�S H�T$pH�L$ H�
H��$�   H�L$0H�
H��HÐSH��0L��L�D$`L���D$     A��� H��� H)�H��0[ÐH�D$(L� �   Ð��   Ð����������   Ð���������H�D$(H�T$0L� H�D$@H��   Ð����H�D$(M)�I9�IF��H��(��N	 ������H��(�H��H��t�*���Y �����H��(��N	 �H��(�H��H��t����Y �������������1�Ð������������AUATUWVSH��8H��$�   L��$�   �H��L��L��L9�D$,�|   M9�swL�l$,�-H���tzH��u
1�f��   �T$,H�H��H9߉U vHI9�vCI��M��H��I)�H����%��H���u��   H��$�   H�H��$�   H�2H��8[^_]A\A]Ð1�H9�����fD  �   �Ő��������AWAVAUATUWVSH��8�H��$�   H��$�   M��I��L�ƉD$$�GM	 L��H)�H�H��H��H��H)�H)�H����   H9���   I9���   L�|$$L�l$+�5H��H)�H9���   H��I��L�������D$$H��H�I9�A�vLH9�vG�M��L���0��H���H��u��   H��$�   H�2H��$�   H�H��8[^_]A\A]A^A_�@ 1�I9�����fD  I9�v;L�|$$�@ �T$$H��H�I9�A�v�M��H���0��H���u���    1�끸   �w�����AUATUWVSH��81�H��$�   �H��I��L��L�ωD$,t_M9�sZL�l$,�6f.�     H����u
�   �   �L$,H��H��H9�       �A�$v"H��tI��H��1�I)�M���#��H�PH��w���H��8[^_]A\A]Ð�������H��(H��L����������������	�H��(Ð������������AWAVAUATUWVSH��HH�|$?L��I��E1�H��L��H�|$(I���?� E1�I��H��H��$�   I���&� I�n�I��H��L��L�`�L�I��6H������H��H��
���H�H9�uI9�t*H9�txI9��   H��H��I��H��L���)�������t�������A�G���~$������A�F���~%��H��H[^_]A\A]A^A_�f�H�T$(I�O���� ��H�T$(I�N��� �˿�����f�     �   �H�T$(I�N�H���� H����������������������H��L��M��������AWAVAUATUWVSH��HH�D$?H��L��1�I��I��H�D$ 1�L��I���� E1�M��H��H�H����� L�x�H)�I��H�D$(H�H��I���Q H��L���Hf�H�H��L�h�M�eL;`�w�@���~L��H���� H�H�P�� H��@�    L�`�B�D( I��I��H��L���)���H9�w(H�XH���HQ H���pQ I��I��H��L��H�������I��H��H���� H���&���H�I9��Z���H���Q H�L$(H�T$ H���?� H��H��H[^_]A\A]A^A_�H��H�H�T$ H���� H���?��H���S H���P �Y H���U H�L$(H�T$ H����� �H����R ��H���ܐ�������������L�9   H�H�@ L9�u�(   �     H���������������H�H�`���������1�L9�sf�     �
��H���I9�u�Ð�������������SH�� H�H���PH��H�� [Ð�       ��������H��(H��L��虾������������	�H��(Ð������������AWAVAUATUWVSH��HH�|$?L��I��E1�H��L��H�|$(I����? E1�I��H��H��$�   I����? I��I�F�L��L��I�,FI�G�M�$G�4H�������H��H�C����H9�H�4FuI9�t&H9�ttI9�tH��H��I��H��L���)�������t�������A�G���~$������A�F���~%��H��H[^_]A\A]A^A_�f�H�T$(I�O���B ��H�T$(I�N���B �˿�����f�     �   �H�T$(I�N�H����B H��� ������������������H��L��M��������AWAVAUATUWVSH��HH�D$?I��L��1�I��I��H�D$ 1�L��H����= E1�I��H��I�$H���> H��H�D$(H�@�H)�L�4FH��������?H9��f  H�?�N I��������?H��H���ND  I�$H��H�p�H��H;p�w�@���~H��L����S I�$1�E1�H�P�f�P�@�    H�p�fD�pI��I��H��L������H9�w2H�xH���eM L9���   H�?�M I��I��H��L��H�������I��H��L���QE H������H�CI9��L���H���M H�L$(H�T$ H���AA L��H��H[^_]A\A]A^A_�H��I�$H�T$ H���A H���P��H���O H����L �U H���#Q H�L$(H�T$ H����@ �H����N ���_V H�����UV �����L�9   H�H�@ L9�u�(   �     H���������������H�H�`���������1�L9�sf�     �
��H���I9�w�Ð�������������SH�� H�H���PH��H�� [Ð���������       AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`�po��D�~H��A��JA��@tA���   �
   E�|$x�H�L$p@��H����@ ����	  �|$h�H�L$`@��H����@ �A����  @8��j  D�t$xH�L$pA���u	H���@	  �Cn�S D8��D$^t
D8so�A	  ��u]D8sHtgH�L$pH�AH;A�;
  H��H�AH�|$p�D$x����H�T$`H��貝�������	  �S E1�1���   f.�     D8sIu�f.�     1�E1�A�����A��D����t
D8sI�E  D8sH�7  D8sr��  E���$  D8spt
D8sq��  �����������  E1�E1��   H�L$pH�AH;A��  H���D$x����H�A1�H�AH9A�C  �|$h�H�L$`@��H����@ �A����  @8��k  �S D�Ǿ   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    ��  �����1�D���   ����E��D$X�  @����  �D$8E1��D$4    �L$@��0�D$]H�|$8
A����  A��/�  D8t$]�
  �AЃ����  �T$49T$X�|  �Չ���9����A��A	�H�L$p�D$4H�AH;A�i  H��H�A�D$@�D$xE1�H�AH9A�  �|$h�H�L$`��H��A��A ���  D8���  L��$�   A�   M���z  E����  @����  H��$0  �     H��$(  �    E��tH��$(  �H��$   foT$pH��$�   H�D$HH��H9�t�H�        H��$   H�ĸ   [^_]A\A]A^A_�A����
��D��t�����A������A��s  H�L$pE1�   H�AH;A������     H�D�D$4�PPH�L$p�D$x����D�D$4H���f����   �l���H�L$pD�t$xH��t
A�����  E���S �����f�     D��1��h���fD  A�F�<	����A�F�<��  �A��������L��$�   E1�M�������L�t$HA��L���'2 H�SM��H�K�7� ����  E��u@��tH��$�    �V���@���M���E����  H��$0  � ����H��$(  �    �?���f�H�L$pA�   H�AH;A�����H��PPH�L$p�D$@H�ɉD$x�����A�   ����1�H�AH9A�M���H�D�D$8�T$4�PH�T$4���D�D$8�*���H�D$`    D������D�t$xH�L$pA��������H�������H�AH;A��  D�0�����     1�H�AH9A����H��PH1҃������H�D$`    D�������A��AA���t����A��e����     H�AH;A�  D�0����f�     A��A������@ @����  H�CrE1��D$4    H�D$@H�D$H�L$_H��H�D$P�C ��t
D8sI�_  D:sH�����L�D$8A��H�L$@�b���H�������H+D$@�P���OT$49T$X�}   �Չ���9����A��A	ωD$4H�L$pH�AH;AsgH���D$x����H�AH�A�D$] H9A��  �|$h�H�L$`��H��A��A �u~:T$]uDL��$�   �����fD  H�L$pE��H�AH;Ar�H��PPH�L$p�D$x����H��u�D�l$]��       �H�L$pD�t$xH�������A��������H�AH;A�V  D�0�����1�H�AH9A�r���H��PH1҃���a���H�D$`    D���P���f�     E��L��$�   �a  H��$�   D�d$]M�fH;D$P�M  H��$�   I9���  �T$]B�0H��$�   L��$�   B�  E1�����1���D���n���H��$�   HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    H�D$8   @ H�L$H�    �a) �]����S �D$^ �   1�E1�E1�������H�D�D$8�T$4�PH�T$4���D�D$8�����H�D$p    �   ����f.�     1�H�AH9A�!���H��PH�������H�D$`    D������1�H�AH9A�����H��PH��������H�D$p    ��������|$4���؀|$^ D�H��$0  ������H��$(  �    ����H�AH;A�1  D�0����fD  �D$^ �&����T$xH���J����S A������H��PH��������H�D$p    A�   �����H�L$HE1�E1�L��H�D$    �?+ H��$�   � ���f�1��   �����ƿ   ����H�D�D$4�PHD�D$4����
  A��������   ����H��PH���A�������H�D$p    H�|$8
������L$@A����������fD  H��PH����D$] �Z���H�D$p    D�l$]�G���H��PP�����H��PH���A���o���H�D$p    �a���H��PH���A���k���H�D$p    D�t$_�W���A��E1�1�L��$�   �D$4    �����A��L��$�   E1�1��D$4    ����E1������H�D$p    E���       ����H��H�D$HH��$�   H��H9�t��? H���]���������������AWAVAUATUWVSH���   �   H��$0  �Ao �Ao	H��$  H���   H��$�   )�$�   )L$p�Mc��D�~H��A��JA��@tA���   �
   E胼$�   �H��$�   @��H����@ ����&	  �|$x�H�L$p@��H����@ �A����  @8��q  D��$�   H��$�   A���u	H���q	  �Cn�S D8��D$dt
D8so�r	  ��u^D8sHthH��$�   H�AH;A�|
  H��H�AǄ$�   ����H�T$pH��$�   H���z��������*	  �S E1�1���   f�D8sIu�f.�     1�E1�A�����A��D����t
D8sI�E  D8sH�  D8sr��  E����  D8spt
D8sq�4	  ����������-	  E1�E1��   H��$�   H�AH;A��  Ǆ$�   ����H��H�A1�H�AH9A�=  �|$x�H�L$p@��H����@ �A����  @8��9  �S D�Ǿ   H�D$@   ��tHc�H�D$@H��$�   ��HǄ$�       H�D$XH��$�   H��$�   Ƅ$�    ��  �D$d1�D���   ������D$L��E��D$H�0  @���(	  �D$@E1��D$<    ��0�D$PH�|$@
A����  A��/��  D8t$P��  �AЃ����  �T$<9T$H�Q  �L$L��)�9����A��A	ωD$<H��$�   H�AH;A�`  Ǆ$�   ����H��H�AE1�H�AH9A�!  �|$x�H�L$p��H��A��A ���  D8��j  L��$�   A�   M���7  E���q  @����       g  H��$@  �     H��$8  �    E��tH��$8  �H��$  fo�$�   H��$�   H�D$XH��H9�t��; H��$  H���   [^_]A\A]A^A_�D  A����
��D��Y�����A������A��x  E1�   �e���H��$�   D��$�   H��t
A�����  E���S �����D��1�����D  A�F�<	�I���A�F�<��  �A�����=���L��$�   E1�M�������L�t$XA��L���'& H�SM��H�K�7� ���/  E��u@��tH��$�    �����@�������E����  �D$dH��$@  ������H��$8  �    �z���f.�     A�   ����D  H�D�D$<�PPH��$�   Ǆ$�   ����D�D$<H���V����   �\���f�     1�H�AH9A�c���H�D�D$@�T$<�PH�T$<���D�D$@�@���H�D$p    D���/���D��$�   H��$�   A��������H�������H�AH;A��  D�0����f�1�H�AH9A�A���H��PH1҃���0���H�D$p    D������A��AA���T����A������     H�AH;A�j  D�0�����f�     H��PPH��$�   Ǆ$�   ����H�������A�   ���� A��A�������@ @���  H�CrE1��D$<    H�D$PH�D$XH��H�D$h�C ��t
D8sI�C  D:sH�����L�D$@A��H�L$P����H�������H+D$P�P���OT$<9T$H��   �L$L��)�9����A��A	ωD$<H��$�   H�AH;A�R  Ǆ$�   ����H��H�AH�A��       D$c H9A��  �|$x�H�L$p��H��A��A �ua:T$cuL��$�   ����E���f�     H��$�   D��$�   H������A��������H�AH;A��  D�0�����fD  1�H�AH9Ar�H��PH1҃��u�H�D$p    D���u���fD  E��L��$�   ��  H��$�   D�d$cM�fH;D$h��  H��$�   I9��  �T$cB�0H��$�   L��$�   B�  E1�����1���D���t���H��$�   HǄ$�       H�D$XH��$�   H��$�   Ƅ$�    H�D$@   @ H�L$X�    �1 �c����S �D$d �   1�E1�E1�������H�D�D$@�T$<�PH�T$<���D�D$@�����HǄ$�       �   �����    1�H�AH9A����H��PH�������H�D$p    D�������1�H�AH9A�����H��PH��������HǄ$�       ������H��PPH��$�   Ǆ$�   ����H�������D�l$c����f��|$<���؀|$d D�H��$@  ������H��$8  �    ����H�AH;A�D  D�0�x���fD  �D$d �������$�   H�������S A�������H��PH��������HǄ$�       A�   ����D  H�L$XE1�E1�L��H�D$    �� H��$�   ������    1��   �L����ƿ   �N���H�D�D$<�PHD�D$<����  A���j����   �q���H��PH���A�������H�|$@
HǄ$�       �v��������A������N���f�H��PH����D$c �B���HǄ$�       D�l$c�,���H��PP����H��PH���A��       ��+���HǄ$�       ����H��PH���A���A���HǄ$�       A������*���A��E1�1�L��$�   �D$<    ����A��L��$�   E1�1��D$<    �}���E1���s���HǄ$�       E���K���H��H�D$XH��$�   H��H9�t�y3 H��������AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`��V��D�~H��A��JA��@tA���   �
   E�|$x�H�L$p@��H����@ ����	  �|$h�H�L$`@��H����@ �A����  @8��j  D�t$xH�L$pA���u	H���@	  �Cn�S D8��D$^t
D8so�A	  ��u]D8sHtgH�L$pH�AH;A�;
  H��H�AH�|$p�D$x����H�T$`H���"��������	  �S E1�1���   f.�     D8sIu�f.�     1�E1�A�����A��D����t
D8sI�E  D8sH�7  D8sr��  E���$  D8spt
D8sq��  �����������  E1�E1��   H�L$pH�AH;A��  H���D$x����H�A1�H�AH9A�C  �|$h�H�L$`@��H����@ �A����  @8��k  �S D�Ǿ   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    ��  �����1�D���   ����E��D$X�  @����  �D$8E1��D$4    �L$@��0�D$]H�|$8
A����  A��/�  D8t$]�
  �AЃ����  �T$49T$X�|  �Չ���9����A��A	�H�L$p�D$4H�AH;A�i  H��H�A�       �D$@�D$xE1�H�AH9A�  �|$h�H�L$`��H��A��A ���  D8���  L��$�   A�   M���z  E����  @����  H��$0  �     H��$(  �    E��tH��$(  �H��$   foT$pH��$�   H�D$HH��H9�t�w/ H��$   H�ĸ   [^_]A\A]A^A_�A����
��D��t�����A������A��s  H�L$pE1�   H�AH;A������     H�D�D$4�PPH�L$p�D$x����D�D$4H���f����   �l���H�L$pD�t$xH��t
A�����  E���S �����f�     D��1��h���fD  A�F�<	����A�F�<��  �A��������L��$�   E1�M�������L�t$HA��L��� H�SM��H�K�� ����  E��u@��tH��$�    �V���@���M���E����  H��$0  � ����H��$(  �    �?���f�H�L$pA�   H�AH;A�����H��PPH�L$p�D$@H�ɉD$x�����A�   ����1�H�AH9A�M���H�D�D$8�T$4�PH�T$4���D�D$8�*���H�D$`    D������D�t$xH�L$pA��������H�������H�AH;A��  D�0�����     1�H�AH9A����H��PH1҃������H�D$`    D�������A��AA���t����A��e����     H�AH;A�  D�0����f�     A��A������@ @����  H�CrE1��D$4    H�D$@H�D$H�L$_H��H�D$P�C ��t
D8sI�_  D:sH�����L�D$8A��H�L$@�қ��H�������H+D$@�P���       �OT$49T$X�}   �Չ���9����A��A	ωD$4H�L$pH�AH;AsgH���D$x����H�AH�A�D$] H9A��  �|$h�H�L$`��H��A��A �u~:T$]uDL��$�   �����fD  H�L$pE��H�AH;Ar�H��PPH�L$p�D$x����H��u�D�l$]�H�L$pD�t$xH�������A��������H�AH;A�V  D�0�����1�H�AH9A�r���H��PH1҃���a���H�D$`    D���P���f�     E��L��$�   �a  H��$�   D�d$]M�fH;D$P�M  H��$�   I9���  �T$]B�0H��$�   L��$�   B�  E1�����1���D���n���H��$�   HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    H�D$8   @ H�L$H�    �� �]����S �D$^ �   1�E1�E1�������H�D�D$8�T$4�PH�T$4���D�D$8�����H�D$p    �   ����f.�     1�H�AH9A�!���H��PH�������H�D$`    D������1�H�AH9A�����H��PH��������H�D$p    ��������|$4���؀|$^ D�H��$0  ������H��$(  �    ����H�AH;A�1  D�0����fD  �D$^ �&����T$xH���|���S A������H��PH��������H�D$p    A�   �����H�L$HE1�E1�L��H�D$    � H��$�   � ���f�1��   �����ƿ   ����H�D�D$4�PHD�D$4����
  A��������   ����H��PH���A�������H�D$p    H�|$8
������L$@A����������fD  H��PH���       ��D$] �Z���H�D$p    D�l$]�G���H��PP�����H��PH���A���o���H�D$p    �a���H��PH���A���k���H�D$p    D�t$_�W���A��E1�1�L��$�   �D$4    �����A��L��$�   E1�1��D$4    ����E1������H�D$p    E������H��H�D$HH��$�   H��H9�t�e' H��������������������AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`��J��D�~H��A��JA��@tA���   �
   E�|$x�H�L$p@��H����@ ����/	  �|$h�H�L$`@��H����@ �A����  @8��z  D�t$xH�L$pA���u	H���Q	  �Cn�S D8��D$Wt
D8so�Q	  ��u]D8sHtgH�L$pH�AH;A�K
  H��H�AH�|$p�D$x����H�T$`H���y�������	  �S E1�1���   f.�     D8sIu�f.�     1�E1�A�����A��D����t
D8sI�U  D8sH�7  D8sr��  E���$  D8spt
D8sq�	  �����������  E1�E1��   H�L$pH�AH;A��  H���D$x����H�A1�H�AH9A�S  �|$h�H�L$`@��H����@ �A����  @8��n  �S D�Ǿ   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    ��  ���  D���   ���E��D$P�"  @���	  �D$8E1�E1�fD�\$T��0�D$@�H�|$8
A���   A��/�  D8t$@�  �AЃ���  �T$Tf9T$P� �        ��H�L$pD�º��  )�A9���D�A��A	�f�D$TH�AH;A�b  H���D$x����H�AE1�H�AH9A�
  �|$h�H�L$`��H��A��A ���  D8���  L��$�   A�   M���s  E����  @����  H��$0  1�f�H��$(  �    E��tH��$(  �H��$   foT$pH��$�   H�D$HH��H9�t�Q# H��$   H�ĸ   [^_]A\A]A^A_�D  A����
��D��i�����A������A��h  H�L$pE1�   H�AH;A�z���H�D�D$T�PPH�L$p�D$x����D�D$TH���c����   �i���H�L$pD�t$xH��t
A�����  E���S �����fD  D��1��h���fD  A�F�<	�	���A�F�<��  �A���������L��$�   E1�M�������L�t$HA��L���w H�SM��H�K�� ����  E��u@��tH��$�    �]���@���T���E����  H��$0  �����f�H��$(  �    �C���H�L$pA�   H�AH;A�����H��PPH�L$p�D$x����H�������A�   ����1�H�AH9A�M���H�D�D$8�T$T�PH�T$T���D�D$8�*���H�D$`    D������D�t$xH�L$pA��������H�������H�AH;A��  D�0�����     1�H�AH9A�%���H��PH1҃������H�D$`    D������A��AA���t����A��`����     H�AH;A�*  D�0����f�     A��A������@ @����  H�CrE1�E1�H�D$@H�D$HfD�T$TH��H�D$X�C ��t
D8sI�       �r  D:sH�����L�D$8A��H�L$@赏��H�������H+D$@�P���O��T$Tf9T$P��   �չ��  )�D��A9����A��A	�f�D$TH�L$pH�AH;AsoH���D$x����H�AH�A�D$V H9A��  �|$h�H�L$`��H��A��A ���   :T$VuHL��$�   �����f.�     H�L$pE��H�AH;Ar�H��PPH�L$p�D$x����H��u�D�l$V�H�L$pD�t$xH�������A��������H�AH;A�V  D�0����1�H�AH9A�n���H��PH1҃���]���H�D$`    D���L���f�     E��L��$�   �c  H��$�   D�d$VM�fH;D$X�M  H��$�   I9���  �T$VB�0H��$�   L��$�   B�  E1�����1���D���^���H��$�   HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    H�D$8   @ H�L$H�    � �M����S �D$W �   1�E1�E1�������H�D�D$8�T$T�PH�T$T���D�D$8�����H�D$p    �   �w���f.�     1�H�AH9A����H��PH�������H�D$`    D�������1�H�AH9A�����H��PH��������H�D$p    ��������|$T���؀|$W D�H��$0  f�����H��$(  �    ����H�AH;A�0  D�0����D  �D$W �����T$xH���p���S A�������H��PH��������H�D$p    A�   �����H�L$HE1�E1�L��H�D$    � H��$�   � ���f�1��   �v����ƿ   �x���H�D�D$T�PHD�D$T����  A��������   ��       ����H��PH���A�������H�D$p    H�|$8
����������A���������D  H��PH����D$V �R���H�D$p    D�l$V�?���H��PP����H��PH���A���_���H�D$p    �Q���H��PH���A���X���H�D$p    A������D���E1�A��L��$�   1�E1�fD�D$T�����E1�A��L��$�   1�fD�L$TE1�����E1������H�D$p    E������H��H�D$HH��$�   H��H9�t�3 H�����������������AWAVAUATUWVSH���   A�   H��$@  �Ao �Ao	H��$   H���   H��$�   )�$�   )�$�   �>��D�{H��A��JA��@tA��A�   �
   DE胼$�   �H��$�   ��H���� ؉���	  ��$�   �H��$�   @��H����@ ����=	  @8���  ��$�   H��$�   ���u	H����	  �Fn�V 8��D$wt	8^o��	  ��u^8^HtdH��$�   H�AH;A��
  H��H�AH��$�   Ǆ$�   ����H��$�   H���l��������	  �V E1�1���   8^Iu�fD  1�E1�A�����A��D����t	8^I��  8^H�Y  8^r��  E���G  8^pt	8^q��	  A�����������	  E1�E1�A�   H��$�   H�AH;A��  Ǆ$�   ����H��H�A1�H�AH9A��  ��$�   �H��$�   @��H����@ �A����  @8���  �V D�ſ   H�D$@   A��tIc�H�D$@H��$�   ��HǄ$�       H�D$hH��$�   H��$�   Ƅ$�    ��  H�       ��|$w H��������D���       �   HE�Ic�H��H�T$P1�H�D$XH��E��H�D$H�}  @���{	  �D$@E1�A�����H�D$8    ��0�D$`fD  H�|$@
����  ��/��  8\$`��  �AЃ����  H�T$8H9T$H��  H�T$PH�H�L$XH)�H9���H�A��A	�H�D$8H��$�   H�AH;A��  H��D��$�   H�AE1�H�AH9A�j  ��$�   �H��$�   ��H���� ���  D8���  H��$�   A�   H���K  E����  @���{  H��$P  H�     H��$H  �    E��tH��$H  �H��$   fo�$�   H��$�   H�D$hH��H9�t�� H��$   H���   [^_]A\A]A^A_�f.�     A��A��
��D�������A��A����A���  E1�A�   �����     H��$�   ��$�   H��t	����#  E���V �����fD  D��1��Q���fD  �C�<	�'����C�<��  �A��������H��$�   E1�H�������H�\$hA��H��� H�VI��H�N�)� ���U  E��u@��tH��$�    �����@���|���E���  H�       ��|$w H��������H��$P  HD�H�H��$H  �    �U���f.�     A�   ����D  H�D�D$8�PPH��$�   Ǆ$�   ����D�D$8H��������   �����f�     1�H�AH9A����H�D�D$@�T$8�PH�T$8���D�D$@�����HǄ$�       D�������f�     ��$�   H��$�   ��������H������H�AH;A�  ��i���f�     �       1�H�AH9A����H��PH1҃�������HǄ$�       ���������A���2����A��=����     H�AH;A�z  ������f.�     H��PPH��$�   D��$�   H���Z���A�   �`���fD  A��A���{���@ @���  H�D$8    H�FrE1�H�D$`H�D$hH��H�D$x�F ��t	8^I�C  :^H�|���L�D$@��H�L$`����H���a���H+D$`�P���O�H�T$8H9T$H��   H�T$PH�H�L$XH)�H9���H�A��A	�H�D$8H��$�   H�AH;A�J  Ǆ$�   ����H��H�AE1�H�AH9A��  ��$�   �H��$�   ��H���� �uUD8�uH��$�   �u��� E���H��$�   ��$�   H���������������H�AH;A��  ������@ 1�H�AH9Ar�H��PH1҃��u�HǄ$�       ������@ E��H��$�   ��  H��$�   E��H;D$xL�c��  H��$�   I9��$  D�<H��$�   L��$�   B�  E1������1�A��D������H��$�   HǄ$�       H�D$hH��$�   H��$�   Ƅ$�    H�D$@   f.�     H�L$h�    �� ������V �D$w �   1�E1�1�����f�H�D�D$@�T$8�PH�T$8���D�D$@�-���HǄ$�       �   �����    1�H�AH9A�����H��PH��������HǄ$�       ������1�H�AH9A�\���H��PH����M���HǄ$�       ���:���H��PPH��$�   Ǆ$�   ����H�������E������f�H�|$8H��H�؀|$w HD�H��$�       P  H��g���H��$H  �    ����f�     H�AH;A�@  �����f.�     �D$w �v�����$�   H���c���V ���\���H��PH��������HǄ$�       A�   �p���fD  H�L$hE1�E1�H��H�D$    �� H��$�   �����    1��   ������ǽ   �����H�D�D$8�PHD�D$8����  ���4����   �`���H��PH������L���H�|$@
HǄ$�       �F���D�������"����    H��PH����?���HǄ$�       E���+���H��PP����H��PH����������HǄ$�       ����H��PH������;���HǄ$�       ������%���A��E1�1�H��$�   H�D$8    �]���A��H��$�   E1�1�H�D$8    �?���E1����5���HǄ$�       D������H��H�D$hH��$�   H��H9�t�A H���������������AWAVAUATUWVSH���   A�   H��$0  �Ao �Ao	H��$  H���   H��$�   )�$�   )L$p�1��D�{H��A��JA��@tA��A�   �
   DE胼$�   �H��$�   ��H���� ؉��	  �|$x�H�L$p@��H����@ �����  @8��a  ��$�   H��$�   ���u	H���p	  �Fn�V 8��D$nt	8^o�v	  ��ub8^HtbH��$�   H�AH;A�z
  H��H�AǄ$�   ����H�T$pH��$�   H����_�������/	  �V E1�1���   �    8^Iu�1�E1�A�����A��D����t	8^I�:  8^H�$  8^r��  E���  8^pt	8^q�D	  A���       ��������<	  E1�E1�A�   H��$�   H�AH;A��  Ǆ$�   ����H��H�A1�H�AH9A�;  �|$x�H�L$p@��H����@ �A����  @8��R  �V D�ſ   H�D$8   A��tIc�H�D$8H��$�   ��HǄ$�       H�D$XH��$�   H��$�   Ƅ$�    ��  D���   Ic�I������1�H��H�D$HL��H��H�D$@E���&  @���$	  �D$8E1�H�D$0    ��0�D$PD  H�|$8
����  ��/��  8\$P��  �AЃ����  H�T$0H9T$@�R  H�T$HH�H��H��H9���H�A��A	�H�D$0H��$�   H�AH;A�I  H��D��$�   H�AE1�H�AH9A�  �|$x�H�L$p��H���� ���  D8��h  H��$�   A�   H���C  E���}  @���s  H��$@  H�     H��$8  �    E��tH��$8  �H��$  fo�$�   H��$�   H�D$XH��H9�t�
 H��$  H���   [^_]A\A]A^A_�f�A��A��
��D��J�����A��A����A��f  E1�A�   �T����     H��$�   ��$�   H��t	�����  E���V �����fD  D��1�����fD  �C�<	�7����C�<��  �A�����,���H��$�   E1�H�������H�\$XA��H���i� H�VI��H�N�y� ���  E��u@��tH��$�    �����@�������E����  H��$@  H� ����H��$8  �    �v��� A�   �����D  H�D�D$0�PPH��$�   Ǆ$�   ����D�D$0H��       �H����   �N���f�     1�H�AH9A�U���H�D�D$8�T$0�PH�T$0���D�D$8�2���H�D$p    D���!�����$�   H��$�   ��������H�������H�AH;A�   �����D  1�H�AH9A�C���H��PH1҃���2���H�D$p    ���"�����A���e����A�����H�AH;A�u  �����D  H��PPH��$�   D��$�   H�������A�   ����fD  A��A�������@ @���  H�FrE1�D�t$oH�D$PH�D$XH�D$0    H��H�D$`�F ��t	8^I�>  :^H�����L�D$8��H�L$P�sv��H�������H+D$P�P���O�H�T$0H9T$@��   H�T$HH�H��H��H9���H�A��A	�H�D$0H��$�   H�AH;A�E  Ǆ$�   ����H��H�AE1�H�AH9A��  �|$x�H�L$p��H���� �uXD8�uH��$�   �����fD  E���H��$�   ��$�   H��������������H�AH;A��  ������@ 1�H�AH9Ar�H��PH1҃��u�H�D$p    �������    E��H��$�   ��  H��$�   E��H;D$`L�c��  H��$�   I9��$  D�4H��$�   L��$�   B�  E1������1�A��D���}���H��$�   HǄ$�       H�D$XH��$�   H��$�   Ƅ$�    H�D$8   f.�     H�L$X�    �� �f����V �D$n �   1�E1�1������f�H�D�D$8�T$0�PH�T$0���D�D$8�����HǄ$�       �   �����    1�H�AH9A�*���H��PH�������H      �D$p    �������1�H�AH9A�����H��PH��������HǄ$�       ������H��PPH��$�   Ǆ$�   ����H�������E������@ H�|$0H��H�؀|$n HD�H��$@  H�����H��$8  �    �����f�     H�AH;A�@  ��z���f.�     �D$n �������$�   H���7W���V �������H��PH��������HǄ$�       A�   ����fD  H�L$XE1�E1�H��H�D$    �$� H��$�   �����    1��   �>����ǽ   �A���H�D�D$0�PHD�D$0����  ���t����   �`���H��PH����������H�|$8
HǄ$�       �����D�������b����    H��PH����B���HǄ$�       E���.���H��PP����H��PH������1���HǄ$�       � ���H��PH������@���HǄ$�       �\$o�*���A��E1�1�H��$�   H�D$0    ����A��H��$�   E1�1�H�D$0    ����E1����}���HǄ$�       D���\���H��H�D$XH��$�   H��H9�t�� H���9������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`�5%��D�kH��A��JA��@��  A��A�
   �  H�D$pH�T$`H��H�D$ H�T$0�T��������  �T$xH�L$ ��T���Vn��8��V �D$Wt	8Fo��  ����  8FH��  H�L$pE1�1���( H�T$0�D$x����H�L$ �S��������  H�D$(   A��tIc�H�D$(H��$�   1�1�I��H      �D$H�t �~  H��$�   ��  �����1҉�A��D$<���   ���D$V��  E1�@����  �D$(E1�L$P��0�D$@H�|$(
����  ��/��  8\$@��  ��0�����  D9l$<�r  E���H�L$p��D9���A�A��H�AA	�H;A�`  H��H�A�D$PH�T$0H�L$ �D$x�R�������~  H��$�   H�y� ��  E����  @����  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�~w H��$�   H�Ę   [^_]A\A]A^A_�f�8FI�����    E1�1��t	8^I�.  8^H�%  8^r��   @���  8^pt	8^q�  A����E�������  E1�1�A�   H�L$pH�AH;A��   H���D$x����H�A1�H�AH9A�3  �|$h�H�L$`@��H����@ �A����  @8���   �   ����H�D$pA�   H�T$`H��H�D$ H�T$0�Q�����������1�E1�1��D$W H�D$(   A�   �[��� ��A��
��@��
���E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$p�D$x����H�������   ����f.�     H�L$p�\$xH��t	����i  @����  �V �L����    �SЀ�	�+����S����  ��W�������H��$�   1�H�y� �|���L��$�   A��L���S� H�VM��H�N胩 ����  E��H��$�   u@��tH�y� �E���@���<���E����  H��$  � ����H��$  �          �.���f.�     H�L$pA�   H�AH;A�����H��PP����1�H�AH9A�����H��T$(�PH�T$(��������H�D$`    D������� �T$xH�L$ �P�����������A���������7������    H�AH;A�:  �����f.�     A����� ���D  1��
���f�     @���  H�FrE1�E1�L$PH�D$@H��$�   H�D$X�F ��t	8^I��   :^H�Q�����H�\$@L�D$(H����j��H���3���H)؍P���O�D9l$<��   E�����D9���A�A��A	�H�L$pH�AH;AswH��H�A�D$PH�T$0H�L$ �D$x��M�������J����T$xH�L$ ��N�����F ���V���8^I�M���E���?  H�L$XA���� H�L$pE1�H�AH;Ar�H��PP�f�D�|$V�e���D  A�   �5���D  H��$�   �    �n� �����f�     1�E1�1��D$W ����H��T$(�PH�T$(��������H�D$p    �   ����@ D���؀|$W DE�H��$  D�(����f�H��$  �    �����T$xH�L$ �M���V �������@ 1��   �����ǽ   ����H��PH���t+���=�����E1�1��������E1�E1�1������1ۉ������H�D$p    ���������H��H��$�   H�T$HH�H��q H��������������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`���D�kH��A��JA��@�   A��A�
   �  H�D$pH�T$`H��H�D$(H�T$8�K�������*  �T      $xH�L$(�|L���Vn��8��V �D$Xt	8Fo�   ����  8FH��  H�L$pE1�1��@  H�T$8�D$x����H�L$(�)K�������2  H�D$0   A��tIc�H�D$0H��$�   1�1�I��H�D$P�/l �~  H��$�   �_  �D$X1�D�d$\D���   ������D$HA��E���D$@�D$L��  @���6  �D$0A��E1��0�D$LH�|$0
���@  ��/�[  8\$L�Q  ��0����E  D9l$@��  �T$HE��H�L$p)�D9���A�A��H�AA	�H;A��  H��H�AH�T$8�D$x����H�L$(�
J��������  H��$�   H�y� ��  E���'  @���  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$PfoT$p��n H��$�   H�Ę   [^_]A\A]A^A_�@ 8FI�����    E1�1��t	8^I��  8^H��  8^r�P  @���s  8^pt	8^q�U  A����E������L  E1�1�A�   H�L$pH�AH;A�R  H���D$x����H�A1�H�AH9A��  �|$h�H�L$`@��H����@ �A���V  @8��9  �   ����H�D$pA�   H�T$`H��H�D$(H�T$8�}H�����������H��$�   1�1�I��H�D$P�i �n H��$�   @����  ���   �D$X @����  H�D$0   1�E1��D$L����D$H����D$\   f.�     @���a  H��$�   E1�E1�H�D$@�F L�fr��t	8^I��   :^H��  L�D$0��L���Vd��H����  L)��P���O�D;l$L��  �T$HD      �l$\)�D9���A�A��A	�H�L$pH�AH;AswH��H�AH�T$8�D$x����H�L$(�LG�������B����T$xH�L$(�4H�����F ���W���8^I�N���E����  H�L$@A���v H�L$pE1�H�AH;Ar�H��PP뉃�A��
��@������E��@��A����@���  H�L$pE1�A�   H�AH;A�����fD  H��PPH�L$p�D$x����H��������   ����f.�     H�L$p�\$xH��t	����i  @����  �V ������    �SЀ�	������S����  ��W��������H��$�   1�H�y� ����L��$�   A��L���c~ H�VM��H�N蓟 ����  E��H��$�   u@��tH�y� �����@�������E����  �D$XH��$  ������H��$  �    �����f�H�L$pA�   H�AH;A�>���H��PP�;���1�H�AH9A�����H��T$0�PH�T$0��������H�D$`    D���q��� �T$xH�L$(�F�����|�����A���������7�����    H�AH;A�*  �����f.�     A���������D  1�����f�     A�   �+���D  A�   �������1�E1��D$X H�D$0   1�H��$�   �    �z �����    1�E1�1��D$X �?���H��T$0�PH�T$0����e���H�D$p    �   �R���@ D���؀|$X DE�H��$  D�(�D���f�H��$  �    �����T$xH�L$(��D���V ���t���@ 1��   �����ǽ   ����H��PH���t/���M�����E1�E1�E1���      ����E1�E1�1�����1ۉ��~���H�D$p    �����������E1�1��_���H��H��$�   H�T$PH�H��h H���η����������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`����D�kH��A��JA��@��  A��A�
   �  H�D$pH�T$`H��H�D$ H�T$0�B��������  �T$xH�L$ �C���Vn��8��V �D$Wt	8Fo��  ����  8FH��  H�L$pE1�1��P H�T$0�D$x����H�L$ �9B��������  H�D$(   A��tIc�H�D$(H��$�   1�1�I��H�D$H�?c �~  H��$�   ��  �����1҉�A��D$<���   ���D$V��  E1�@����  �D$(E1�L$P��0�D$@H�|$(
����  ��/��  8\$@��  ��0�����  D9l$<�r  E���H�L$p��D9���A�A��H�AA	�H;A�`  H��H�A�D$PH�T$0H�L$ �D$x�(A�������~  H��$�   H�y� ��  E����  @����  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�f H��$�   H�Ę   [^_]A\A]A^A_�f�8FI�����    E1�1��t	8^I�.  8^H�%  8^r��   @���  8^pt	8^q�  A����E�������  E1�1�A�   H�L$pH�AH;A��   H���D$x����H�A1�H�AH9A�3  �|$h�H�L$`@��H����@ �A����  @8���   �   ����H�D$pA�   H�T$`H��H�D$ H�T$0�      ?�����������1�E1�1��D$W H�D$(   A�   �[��� ��A��
��@��
���E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$p�D$x����H�������   ����f.�     H�L$p�\$xH��t	����i  @����  �V �L����    �SЀ�	�+����S����  ��W�������H��$�   1�H�y� �|���L��$�   A��L����v H�VM��H�N�� ����  E��H��$�   u@��tH�y� �E���@���<���E����  H��$  � ����H��$  �    �.���f.�     H�L$pA�   H�AH;A�����H��PP����1�H�AH9A�����H��T$(�PH�T$(��������H�D$`    D������� �T$xH�L$ �>�����������A���������7������    H�AH;A�:  �����f.�     A����� ���D  1��
���f�     @���  H�FrE1�E1�L$PH�D$@H��$�   H�D$X�F ��t	8^I��   :^H�Q�����H�\$@L�D$(H���xY��H���3���H)؍P���O�D9l$<��   E�����D9���A�A��A	�H�L$pH�AH;AswH��H�A�D$PH�T$0H�L$ �D$x�r<�������J����T$xH�L$ �Z=�����F ���V���8^I�M���E���?  H�L$XA���t H�L$pE1�H�AH;Ar�H��PP�f�D�|$V�e���D  A�   �5���D  H��$�   �    ��q �����f�     1�E1�1��D$W ����H��T$(�PH�T$(�������      �H�D$p    �   ����@ D���؀|$W DE�H��$  D�(����f�H��$  �    �����T$xH�L$ �O<���V �������@ 1��   �����ǽ   ����H��PH���t+���=�����E1�1��������E1�E1�1������1ۉ������H�D$p    ���������H��H��$�   H�T$HH�H��&` H���N�����������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`�E��D�kH��A��JA��@��  A��A�
   �  H�D$pH�T$`H��H�D$(H�T$8�$:��������  �T$xH�L$(�;���Vn��8��V �D$Wt	8Fo��  ����  8FH��  H�L$pE1�1��� H�T$8�D$x����H�L$(�9��������  H�D$0   A��tIc�H�D$0H��$�   1�1�I��H�D$H�Z �~  H��$�   ��  ���  �A���D$P���   ���D$V��  E1�@����  �D$0E1��0�D$@f�H�|$0
����  ��/��  8\$@��  ��0�����  fD9l$P�v  E����  )�A��9�H�L$p��A�A��A	�H�AH;A�^  H��H�AH�T$8�D$x����H�L$(�8�������|  H��$�   H�y� ��  E����  @����  H��$  E1�fD� H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�] H��$�   H�Ę   [^_]A\A]A^A_�8FI����fD  E1�1��t	8^I�.  8^H�%  8^r��   @���  8^pt	8^q�  A����E�������  	      E1�1�A�   H�L$pH�AH;A��   H���D$x����H�A1�H�AH9A�3  �|$h�H�L$`@��H����@ �A����  @8���   �   ����H�D$pA�   H�T$`H��H�D$(H�T$8�7�����������1�E1�1��D$W H�D$0   A�   �[��� ��A��
��@��
���E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$p�D$x����H�������   ����f.�     H�L$p�\$xH��t	����i  @����  �V �L����    �SЀ�	�&����S����  ��W�������H��$�   1�H�y� �~���L��$�   A��L���cn H�VM��H�N蓏 ����  E��H��$�   u@��tH�y� �G���@���>���E����  H��$  �����f�H��$  �    �/����     H�L$pA�   H�AH;A�����H��PP����1�H�AH9A�����H��T$0�PH�T$0��������H�D$`    D������� �T$xH�L$(�6�����������A���������7������    H�AH;A�:  �����f.�     A����� ���D  1��
���f�     @���  H�FrE1�E1�H�D$@H��$�   H�D$X�F ��t	8^I��   :^H�U�����H�\$@L�D$0H����P��H���7���H)؍P���O�fD9l$P��   E����  )�A��9���A�A��A	�H�L$pH�AH;AswH��H�AH�T$8�D$x����H�L$(��3�������I����T$xH�L$(��4�����F ���O���8^I�F���E���< 
       H�L$XA���l H�L$pE1�H�AH;Ar�H��PP�D�|$V�g���@ A�   �5���D  H��$�   �    �~i �����f�     1�E1�1��D$W ����H��T$0�PH�T$0��������H�D$p    �   ����@ D���؀|$W DE�H��$  fD�(�����H��$  �    �����T$xH�L$(��3���V �������@ 1��   �����ǽ   ����H��PH���t+���=�����E1�1��������E1�E1�1������1ۉ������H�D$p    ���������H��H��$�   H�T$HH�H��W H���Φ����������������AWAVAUATUWVSH��   H��$  �Ao �Ao	H��$�   H���   H��$�   )�$�   )L$p����D�sH��A��JA��@��  A��A�
   �b  H�D$pL��$�   H��H�D$0L���1��������  ��$�   L���2���Vn��8��V �D$_t	8Fo�;  ���#  8FH�*  H��$�   E1�1��H H�T$0L��Ǆ$�   �����01��������  fD  H�D$(   A��tIc�H�D$(H��$�   1�1�I��H�D$`�0R �~  H��$�   ��  H�       ��|$_ H��������D���   HE�Ic�H��H�T$@1�H�D$HH��E��H�D$8H�D$P��  @����  �D$(A��E1��0�D$PfD  H�|$(
���A  ��/�\  8\$P�R  ��0����F  L9d$8��  L�d$@H�H�T$HH)�L9���I�A��A	�H��$�   H�AH;A��  H��H�AH�T$0L��Ǆ$�   ������/�������  H��$�   H�y� ��  E��      �  @���  H��$   H�     H��$  �    ��tH��$  �H��$�   H��H�T$`fo�$�   ��T H��$�   H�Ĩ   [^_]A\A]A^A_��    8FI������    1�E1�A��D��D  ��t	8^I��  8^H��  8^r�q  E����  8^pt	8^q��  A�����������  E1�E1�A�   H��$�   H�AH;A�t  Ǆ$�   ����H��H�A1�H�AH9A��  �|$x�H�L$p@��H����@ �A���q  @8��  D�ſ   �;���H�D$pA�   L��$�   H��H�D$0L���8.�����������H��$�   1�1�I��H�D$`�UO �n H��$�   @����  ���   �D$_ @����  H��������1�E1�H�D$(   H�D$PH��������H�D$HH�D$@   fD  @����  H�FrE1�E1�H�D$8H��$�   H�D$h�F ��t	8^I��   :^H�u  ��H�\$8L�D$(H����I��H���W  H)؍P���O�L;d$P��  L�d$@H�H�T$HH)�L9���I�A��A	�H��$�   H�AH;A�f  H��H�AH�T$0L��Ǆ$�   ������,������������$�   L����-�����F ���E���8^I�<���E����  H�L$hA���e E1��{����    A��A��
��D��������A��A����A��  E1�A�   �����     H��$�   ��$�   H��t	�����  E����  �V ������SЀ�	������S����h  ��W��������H��$�   1�H�y� �#���L��$�   A��L���Cd H�VM��H�N      �s� ���K  E��H��$�   u@��tH�y� �����@�������E����  H�       ��|$_ H��������H��$   HD�H�H��$  �    ����A�   �.���D  H�D�D$(�PPH��$�   Ǆ$�   ����D�D$(H���r����   �x���f�     1�H�AH9A����H�D�D$8�T$(�PH�T$(���D�D$8�\���H�D$p    D���K�����$�   L���+�����6���fD  ��A���������7�A���H�AH;A�V  ��C���fD  H��PP�l���D  A��A������@ D��1��&���fD  A�   ����D  A�   �h�����1�E1��D$_ H�D$(   1�H��$�   �    �` �����    1�E1�1��D$_ �����H�D�D$8�T$(�PH�T$(���D�D$8�+���HǄ$�       �   ����fD  H��PP����D  L��H�؀|$_ LE�H��$   L� ������H��$  �    ������$�   L���N*���V ������ 1��   �����ǽ   ����H�D�D$(�PHD�D$(���t/���������E1�E1�E1��$�����E1�E1�1�����1ۉ�����HǄ$�       �����������E1�1������H��H��$�   H�T$`H�H��N H���0�������������������AWAVAUATUWVSH��   H��$  �Ao �Ao	H��$�   H���   H��$�   )�$�   )L$p�"���D�sH��A��JA��@��  A��A�
   �=  H��$�   H�T$pH��H�D$(H�T$8��'��������  ��$�   H�L$(��(���Vn��8��V �D$gt	      8Fo�  ����  8FH�  H��$�   E1�1��� H�T$8Ǆ$�   ����H�L$(�'�������  H�D$0   A��tIc�H�D$0H��$�   1�1�I��H�D$X�H �~  H��$�   �  D���   Ic�H������1�I��H�D$HH��I��H�D$@E����  E1�@����  �D$0E1�A�σ�0�D$`H�|$0
����  ��/��  8\$`��  ��0�����  L9d$@�W  L�d$HH�H��H��L9���I�A��A	�H��$�   H�AH;A��  H��H�AH�T$8D��$�   H�L$(�d&�������z  H��$�   H�y� �`  E����  @����  H��$   H�     H��$  �    ��tH��$  �H��$�   H��H�T$Xfo�$�   �FK H��$�   H�Ĩ   [^_]A\A]A^A_�f.�     8FI������    E1�1��t	8^I�.  8^H�%  8^r��   @���  8^pt	8^q�  A����E������  E1�1�A�   H��$�   H�AH;A��  Ǆ$�   ����H��H�A1�H�AH9A�-  �|$x�H�L$p@��H����@ �A����  @8���   �   �i���f�     H��$�   A�   H�T$pH��H�D$(H�T$8�$�����������1�E1�1��D$g H�D$0   A�   �(������A��
��@������E��@��A����@���  E1�A�   �����     H��$�   ��$�   H��t	�����  @����  �V �v�����SЀ�	�F����S����H  ��W����:���H��$�   1�H�y� �����L��$�   A��L��      �C\ H�VM��H�N�s} ���+  E��H��$�   u@��tH�y� �i���@���`���E����  H��$   H� ����H��$  �    �R���f�     A�   ����D  H��PPH��$�   Ǆ$�   ����H�������   ����@ 1�H�AH9A����H��T$0�PH�T$0��������H�D$p    D��������    ��$�   H�L$(��#����������     ��A���������7�����H�AH;A�V  ��c���fD  H��PP�
���D  A����� ���D  1������f�     @���-  H�FrE1�E1�L$`H�D$PH��$�   H�D$h�F ��t	8^I��   :^H�!�����H�\$PL�D$0H���>��H������H)؍P���O�L9d$@��   L�d$HH�H��H��L9���I�A��A	�H��$�   H�AH;A��   H��H�A�D$`H�T$8H�L$(��$�   �!�������.�����$�   H�L$(�w"�����F ���C���8^I�:���E���<  H�L$hA���Y E1��w����E���n����     A�   ����D  H��$�   �    �.W �����f�     1�E1�1��D$g �~���H��T$0�PH�T$0��������HǄ$�       �   �����H��PP�	���D  L��H�؀|$g LE�H��$   L� �z����H��$  �    �������$�   H�L$(�l!���V �������1��   ������ǽ   �����H��PH���t+��������E1�1��������E1�E1�1������1ۉ�����HǄ$�       ����������H��H��$�   H�T$XH�H��CE H��      �k��������������AWAVAUATUWVSH��xH��$�   �Ao �Ao	H��$�   H���   H�L$f)D$PL�|$@)L$@�f���L�d$PL��L��H���s������  ��1�E1�1�f�H�D$g1�1�I��H�D$8�@ �~  H�D$h��  ���   ���D$/�H  @���  �V H�FrE1�H�D$ H�D$hH�D$0D  ��t	8^I��  8^H�:  H�L$ ��A�
   �w;��H����  H+D$ H��$�   �P0���&W �|$/A��H�L$PH�AH;A�9  H��H�AL��L���D$X����������'  H�\$hH�C�H��tJ@����  E����  L�t$hA��L���V H�\$hH�VM��H�N��w ��uH��$�   �    H��$�   H�K�H�T$8foT$P�`C H��$�   H��x[^_]A\A]A^A_��    @����  E1��C���<	wn��0���tfH��$�   ��0���V �   H�L$PH�AH;A�/  H��H�AL��L���D$X�����|����������T$XL���h���ÍC���<	v�8^H�c  8��   t8��   �����D����@ ������H��$�   �e   �U H�L$PH�AH;A�^  H��H�AL��L���D$X�����������  �T$XL������8Fo���A  8Fn�-   �8  A�������L�t$h�p����H�\$hA�H�C���  H��tH�L$0A����T H��$�   �.   ��T H�L$P�l$/H�AH;A�����H��PP�����fD  �T$XL���D�����V �9���f�     8��   t8��   �����H�\$hD���@ �H�C������H��t	@���6  H��$�   �e   �      TT H�L$P��� L��L���D$X������������  �T$XL������No���V 8�tu8FntpA�������     �+   H��$�   ��S H�L$PA��H�AH;A�����H��PP�����D���  E���  H�L$0A���S E1�E1�����f���t	8FI�3  8FH�z���1�8�H��$�   �T+�rS A���M���f.�     ��D������H��$�   �.   �CS E1��   ����fD  H�L$0A���"S ����H��PP����f�L�t$h�    L���P �N���f�     �T$XL���t���No���V 8���   8Fn��   1�E1�A�������t	8^I��   8^H��   8^r�   @��t:H�L$PA��H�QH;QsWH��H�QL��L��D�t$X������t�ŉ�����f�H��$�   �0   �NR 벋T$XL��   �����V ���r���H��PP��     1��I���f�     ��t	8FI�:���8FH�1���1�8�H��$�   ��1�E1�T+��Q H�L$P�c� L��L���D$X�����P������������T$XL���:���V �������H��$�   E1�1�H��$�   H� L�@��P H�\$hH�{� ����������f�     A�։������fD  H�\$hL�t$hH�{� ���������H�\$hH�C�L�t$hH���n�������H��H�D$hH�T$8H�H���= H������������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P`H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$      PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PPH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PXH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PHH��H��`[ÐSH��`L�$  H��Ao�Ao	L��$�   H�@(H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L�  H��Ao�Ao	L��$�   H�@H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@0H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@ H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@8H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@@H��      )\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u�(���H��H��`[���H��H��`[Ð���UWVSH��   H��$�   I� �AoI�X�n)D$@L�L$@H��L�D$P��ᵃ��NH�L$`H�D$PH�D$xH�D$0H��$�   H�t$ H�\$XH�D$(�����T$hH�    ����H�D$`H!ˉnH�L$xH	�H��$�   H�H��H�_H�
H�Ĉ   [^_]Ð��������������AWAVAUATUWVSH��   H��$   M�QM�M�`M�	I���@L��$�   L��$�   L��$�   L��$�   ��   H��$(  L�L$PH�L$pL��$�   H�D$ L�D$0L�L$PL�D$`L�\$`H�|$(Ǆ$�   ����L�d$hL�T$X����H�D$pH��$�   �D$x��$�   ��$�   ���   H��$0  ��'fo�$�   L��AE H�ĸ   [^_]A\A]A^A_�H���   A�   A�   H��$�   ����A�����H�x@ I��A��H�x0 A��1�E���  ��$�   �H��$�   ��H���� ؉���  ��$�   �H��$�   @��H����@ �����  @8��'  ��$�   H��$�   ���u	H����  E����   I�V8�*8�A���/  E���T  I�V(8*A���     D��D��d  H��$�   H��H�AH;A�
  H��H�AE��D��$�   ��   I9n@A��E����   E��E�������1�E��tI9n@u	H����  E��tI9n0u	H����  H��$0  ��� ��  H��$(  �    �A���@ I�V(�*8�A���<���E����  I9n@�y  H���p  H��$0  �  1�       H��$(  �������A��I9n0A��A���=���E������������1�H�AH9A�p���H�D�L$OD�D$N�PHA�����D�D$N���D�L$O�E���HǄ$�       ���2����1�H�AH9A�����H�D�L$OD�D$N�PHA�����D�D$N���D�L$O�����HǄ$�       ������f�H�AH;A��   � �����f.�     H��$0  H��$�   H��$�   � H��$(  �    �����������H��$(  ������f.�     H��PPA����������E��t*I9n0��   H��$0  �  H��$(  �    ����f�H��$0  �  H��$(  �    �_���f�H�D�L$OD�D$N�PHA�����D�D$N���D�L$O����HǄ$�       �����������   ����H���l���H��$0  � 1������H��$0  E��� t
I9n0�K�����������H��$0  ��鐐�������AWAVAUATUWVSH��   I�8I�pM�!M�qL��$�   H��I��1�1�M����. H��$�   �    H��H��$�   �C H��$  H�L$pH�\$0L��L�L$PH�|$`L�D$`H�t$hL�d$PH�D$(H��$   L�t$XH�D$ �N���H�    ����H�|$p�D$xH!�I��H	��]s L��$  M��H��$�   H��$  H��$�   �Y ���@��H����@ ��D$O��   A�����M��t��uK@8�uH��$  �H��$�   L�} �����H�]��A���~=H��H�Ę   [^_]A\A]A^A_�fD  1�I�T$I9T$r�I�$L���PH������H��L���1 �f�1�H�GH9G�e���H�H���PH�T$O���A�    L      E�D��B���H��H��$�   L��H�H��F1 H���n�����������������AWAVAUATUWVSH��   I�8I�pM�!M�qL��$�   H��I��1�1�M����, H��$�   �    H��H��$�   �A H��$  H�L$pH�\$0L��L�L$PH�|$`L�D$`H�t$hL�d$PH�D$(H��$   L�t$XH�D$ �^���H�    ����H�|$p�D$xH!�I��H	��mq L��$  M��H��$�   H��$  H��$�   �X ���@��H����@ ��D$O��   A�����M��t��uK@8�uH��$  �H��$�   L�} �����H�]��A���~=H��H�Ę   [^_]A\A]A^A_�fD  1�I�T$I9T$r�I�$L���PH������H��L���/ �f�1�H�GH9G�e���H�H���PH�T$O���A�    LE�D��B���H��H��$�   L��H�H��V/ H���~~����������������ATUWVSH��   �Ao �Ao	H��$�   H��$�   H��I��)�$�   1�1�I��)L$p��* H��$�   �    H��H��$�   �? H��$�   H�L$`H�l$0L��fo\$pH�\$(L�L$@fo�$�   L�D$P)\$@H�D$ )T$P�f���H�D$`H��$�   �D$h��$�   �yo H��$   I��I��H��$�   H��$�   ��W H�T$pH��$�   ������t�H��$�   �����fo�$�   '��A���~H��H�Ġ   [^_]A\�f.�     H��H����- ��H��H��$�   H��H�H���- H���}�����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �~���H��H��`[Ð����      SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ 螻��H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �.���H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �N���H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �n���H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ ����H��H��`[Ð����AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`�����D�vH��A��JA��@tA���   �
   E�f�|$x�H�L$p@��H����@ ����
  f�|$h�H�L$`��H���� Љ���	  @8��k	  H�L$pD�l$xH��tfA����L
  ���   �S fD9��D$_tfD9��   �X
  ��uVfD9kHt]H�L$pH�AH;A�Y  H��H�AH�|$p�����H�T$`H��f�t$x�F�������
  �S E1�1���   fD9kJu��    E1�1���tfD9kJ�V  fD9kH�Q  fD9��   ��  @���:  fD9��   tfD9��   ��	  ����E������
  E1�1��   H�L$pH�AH;A��  H��A�����H�AfD�\$xH�AH;A�O  � E1�f����/  f�|$h�H      �L$`��H���� Љ���  A8��h  �S �   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    ��  1Ҹ����D���   ��E���D$X��  @���R	  �D$8�D$^ �D$4    D�x0H�|$8
A���3  fA��/�X  fE9��N  ��0����B  �T$4�L$X9��  �Չ���9����A��L$^�D$4H�L$pH�AH;A��  H��A�����H�AfD�L$xH�AH;A�\  � E1�f����c  f�|$h�H�L$`��H��A��A ��%  A8���  L��$�   A�   H��$�   M����  @���  E���  H��$0  �     H��$(  �    E��tH��$(  �H��$   foT$pH�D$@H��H9�t�:� H��$   H�ĸ   [^_]A\A]A^A_Ã���
��@��R���E��@�ǃ���@���  H�L$pE1�   H�AH;A�j���H��PPH�L$pA�����fD�T$xH���^���A�   �q���H�L$pD�l$xH��tfA����%  @���S ������     1��j���f�     H�AH;A�r  � 1�f����2���H�D$`    ���"��� A�U�f��	�����A�U�f����  ��W���������     L��$�   E1�H��$�   M���W���H�D$@I�mE��H��H9���  H��$�   H9��
  F�<)H��$�   H��$�   L�D$@�( H�SH�K� Z ���K  E��H��$�   u@��tH��$�    �����@��������|$^ ��  H��$0  � ����H��$(  �    ������      H�L$p�D$^H�AH;A����H��PPH�L$pA�����fD�D$xH������A�   ����D�l$xH�L$pfA����d���H���[���H�AH;A��  D�(fA����>���H�D$p    H�|$8
��������  �p���f�H�AH;A�  � 1�f��������H�D$`    D������f�H�AH;A��  D�(fA��������H�D$p    ����D  A��������D  A��AfA��������7����f�     H�D$p    A�   ����@����  H���   �D$^ H�D$HH�D$@�D$4    H��H�D$P�C ����   fD9kJ��   E��L��$�   H��$�   ��  H;L$PM�}�}  H��$�   I9���  F�$)H��$�   E1�L��$�   B�8 H�L$pH�AH;A��   H�������H�Af�T$xH�AH;A��  � E1�f����@  f�|$h�H�L$`��H��A��A ��"  D8���   L��$�   H��$�   �;����fD;kH�����H�D$HH�T$8fD9(tD  H��H�������fD9(u�H+D$H�L$4H���P���O�9L$X��   H�L$pD�t$^H�AH;A�(���H��PPH�L$p�����f�D$xH������E���2���H�L$pD�l$xH���o���fA����d���H�AH;A�b  D�(fA����G���H�D$p    �9���D  �T$4������9����A��L$^�D$4�}���H�AH;A�s  � 1�f��������H�D$`    D������H�L$@E1�E1�L��H�D$    �c� H��$�   �
���1����z���H��$�   HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    H�      D$8   �H�L$@�    豏 �l����S �D$_ �   1�E1�E1�������   ����fD  H��PH����D  H��PH����D  H�AH;A��  � 1�f����#���H�D$`    ������ H�AH;A��  � 1�f��������H�D$p    ������� H�D$p    A�   �����t$4���؀|$_ D�H��$0  ������H��$(  �    ����f.�     H�AH;A�p  D�(fA��������H�D$p    ����D  �D$_ �����T$xH���)����S A�������H�D$p    E������1��   ����H�L$@E1�E1�L��H�D$    �t� H��$�   �����H��PH����H��PH������ƿ   �t���H��PHA���	���H��PH�2���H��PH�����   �t���A��L��$�   1��D$^ H��$�   �D$4    �z���A���D$^ 1�L��$�   H��$�   �D$4    �S���H��PHA������E1����;���H��PP����H��PH�����H��PH�!���H��PHA������H��PHA������H��H�D$@H��$�   H��H9�t膦 H����m����������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`�����D�vH��A��JA��@� 
  A��A�
   ��  H�l$`H�|$pH��H�����������6
  H�L$pD�l$xH��tfA�����
  ���   �S fD9��D$[t
fD9��   uf��uRfD9kHt[H�L$pH�AH;A��  H��H�A�����H��H��f�t$x���������|
  �S 1�1���   @       fD9kJu�f�     1�1���tfD9kJ�(	  fD9kH�r  fD9��   ��  @���[  fD9��   tfD9��   �;
  A����E������q
  1�1�A�   H�L$pH�AH;A��  H��A�����H�AfD�\$xH�AH;A�	  � E1�f����_  f�|$h�H�L$`��H���� Љ���  A8���  �S �   H�D$8   A��tIc�H�D$8H��$�   ��HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    �P  1��|$[ D�d$\��1�����D$PA���    �D$@�D$T�=  @����	  �D$8E1��D$4    ��0f�D$TH�|$8
A���<  fA��/�a  fD;l$T�U  ��0����I  �T$49T$@�  �L$PA��)�9���Ѓ�A	�H�L$p�D$4H�AH;A�  H��A�����H�AfD�L$xH�AH;A��  � E1�f�����  f�|$h�H�L$`��H��A��A ��=  A8���  L��$�   A�   H��$�   M����  D  @���#  ���  H��$0  �     H��$(  �    E��tH��$(  �H��$   foT$pH�D$HH��H9�t�n� H��$   H�ĸ   [^_]A\A]A^A_�f�H�l$`A�   H�|$pH��H���e������L����s H��$�   HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    @����  ���   1�1���D$[��  �t$[1��D$[ E1��D$T����D$P���H�D$8   �D$\   �     @����  H�D$HL���   E1��D$4    H��H�D$@�C ���O  fD9kJ�D  ��L��$�         H��$�   ��  H;L$@M�l$��  H��$�   I9���  B�,!H��$�   1�L��$�   B�( H�L$pH�AH;A�?  H�������H�Af�T$xH�AH;A��  � E1�f�����  f�|$h�H�L$`��H��A��A ��@  A8������H�L$pD�l$xH������fA�������H�AH;A��  D�(fA��������H�D$p    ������     ��A��
��@��2���A��@��E����@���  H�L$p1�A�   H�AH;A�J���H��PPH�L$pA�����fD�T$xH���>���A�   �Q���D�l$xH�L$pfA���u	H���5  @���S �|����     1��J���f�     H�AH;A�"  � 1�f�������H�D$`    ������ A�U�f��	�����A�U�f���  ��W���������     L��$�   E1�H��$�   M���T���H�D$H@�l$8M�t$H��H9���  H��$�   I9��K  B�,!H��$�   L��$�   L�D$HB�0 H�SH�K�,K ����  ��H��$�   u@��tH��$�    �����@�������E���E  1��|$[ H��$0  ������H��$(  �    �����D  H�L$pA�   H�AH;A�����H��PPH�L$pA�����fD�D$xH�������A�   ����H�L$pD�l$xH���L���fA����A���H�AH;A�#  D�(fA����$���H�D$p    H�|$8
��������  �_����H�AH;A�/  � 1�f��������H�D$`    D������f�H�AH;A�!  D�(fA��������H�D$p    ����D        ��������fD  A��AfA��������7����f�     H�D$p    A�   ����fD;kH�����L��H�T$8fD9(t H��H�������fD9(u�L)��L$4H���P���O�9L$TsCH�L$pA�   H�AH;A�����H��PPH�L$p�����f�D$xH�������A�   �������L$P�T$4�T$\)�9���Ѓ�A	ωD$4�_���H�AH;A�  � 1�f��������H�D$`    D������H�L$HE1�E1�L��H�D$    �� H��$�   �����@ A�   ����1�A�������H��$�   HǄ$�       H�D$HH��$�   H��$�   Ƅ$�    H�D$8   H�L$H�    �0� �����S E1�1�1��D$[ �F���fD  �   �V���fD  H��PH�����D  H��PH�����D  H�D$p    A�   �1����t$4���؀|$[ D�H��$0  �����H��$(  �    �V���f.�     H�AH;A�g  D�(fA����-���H�D$p    �����T$xH�������S A������H�D$p    A�   �����1��   �M���H�L$HE1�E1�L��H�D$    �`� H��$�   ����H��PH�����H��PH�E����ƿ   ����H��PHA�������H��PH�r���H��PH������   �3���E1�1�1��D$[ H�D$8   �Z���L��$�   �D$4    E1�1�H��$�   A�   ����A��E1�1�L��$�   H��$�   �D$4    �����H��PHA�������E1�������H��PP�)���H��PHA���*���H��PHA������H��H�D$HH��$�   H��H9�t�o� H����`�      ��������AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`�н��D�vH��A��JA��@tA���   �
   E�f�|$x�H�L$p@��H����@ �����	  f�|$h�H�L$`��H���� Љ���	  @8��;	  H�L$pD�l$xH��tfA����
  ���   �S fD9��D$_tfD9��   �(
  ��uVfD9kHt]H�L$pH�AH;A��
  H��H�AH�|$p�����H�T$`H��f�t$x�V���������	  �S E1�1���   fD9kJu��    E1�1���tfD9kJ�&  fD9kH�a  fD9��   ��  @���J  fD9��   tfD9��   ��	  ����E�������	  E1�1��   H�L$pH�AH;A��  H��A�����H�AfD�\$xH�AH;A�  � E1�f�����  f�|$h�H�L$`��H���� Љ���  A8��x  �S �   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    �P  1Ҹ����D���   ��E���D$X�v  @����  �D$8�D$^ �D$4    D�x0H�|$8
A���C  fA��/�h  fE9��^  ��0����R  �T$4�L$X9���  �Չ���9����A��L$^�D$4H�L$pH�AH;A��  H��A�����H�AfD�L$xH�AH;A�  � E1�f����3  f�|$h�H�L$`��H��A��A ���  A8���  L��$�   A�   M����  D  E����  @����  H��$0  �     H��$(  �    E��tH��$(  �H      ��$   foT$pH��$�   H�D$@H��H9�t�E� H��$   H�ĸ   [^_]A\A]A^A_�f�     ����
��@��D���E��@�ǃ���@��x  H�L$pE1�   H�AH;A�\���H��PPH�L$pA�����fD�T$xH���P���A�   �c���f�H�L$pD�l$xH��tfA�����  @���S ������     1��Z���f�     H�AH;A�2  � 1�f����"���H�D$`    ������ A�U�f��	�����A�U�f����  ��W���������     L��$�   E1�M���L���L�|$@A��L���+ H�SM��H�K�;@ ���F  E��u@��tH��$�    ����@�������|$^ ��  H��$0  � ����H��$(  �    ����@ H�L$p�D$^H�AH;A�C���H��PPH�L$pA�����fD�D$xH���7���A�   �J���D�l$xH�L$pfA��������H�������H�AH;A�u  D�(fA����n���H�D$p    H�|$8
��������  ����f�H�AH;A��  � 1�f��������H�D$`    D�������f�H�AH;A��  D�(fA��������H�D$p    �����D  A���������D  A��AfA���Q�����7�����f�     H�D$p    A�   �����@����  H���   �D$^ H�D$HH�D$@�D$4    H��H�D$P�C ����   fD9kJ��   E��L��$�   �v  H��$�   M�}H;D$P�}  H��$�   I9���  F�$(H��$�   E1�L��$�   B�8 H�L$pH�AH;A��   H�������H�Af�T$xH�A      H;A��  � E1�f����@  f�|$h�H�L$`��H��A��A ��"  D8���   L��$�   �k���f�     fD;kH����H�D$HH�T$8fD9(tD  H��H�������fD9(u�H+D$H�L$4H���P���O�9L$X��   H�L$pD�t$^H�AH;A�(���H��PPH�L$p�����f�D$xH������E���2���H�L$pD�l$xH���o���fA����d���H�AH;A�  D�(fA����G���H�D$p    �9���D  �T$4������9����A��L$^�D$4�}���H�AH;A�J  � 1�f��������H�D$`    D������H�L$@E1�E1�L��H�D$    �y H��$�   �
���1��������H��$�   HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    H�D$8   �H�L$@�    ��u �����S �D$_ �   1�E1�E1��2�����   ����fD  H��PH�����D  H��PH�����D  H�AH;A��  � 1�f����S���H�D$`    ���C��� H�AH;A��  � 1�f�������H�D$p    ������� H�D$p    A�   �����t$4���؀|$_ D�H��$0  �����H��$(  �    ����f.�     H�AH;A�-  D�(fA��������H�D$p    ����D  �D$_ �6����T$xH���i����S A������H�D$p    E������1��   �����H��PH�����H��PH�����ƿ   �����H��PHA���2���H��PH�[���H��PH����A���D$^ 1�L��$�   �D$4    �����H��PHA������A��L��$�   �D      $^ 1��D$4    ����E1�������H��PP����H��PH�o���H��PH�4���H��PHA�������H��PHA�������H��H�D$@H��$�   H��H9�t�	� H���qT���AWAVAUATUWVSH��   �   H��$   �Ao �Ao	H��$   H���   H��$�   )D$p)L$`�p���D�vH��A��JA��@tA���   �
   E�f�|$x�H�L$p@��H����@ �����	  f�|$h�H�L$`��H���� Љ���	  @8��K	  H�L$pD�l$xH��tfA����,
  ���   �S fD9��D$_tfD9��   �8
  ��uVfD9kHt]H�L$pH�AH;A��
  H��H�AH�|$p�����H�T$`H��f�D$x�����������	  �S E1�1���   fD9kJu��    E1�1���tfD9kJ�5  fD9kH�a  fD9��   ��  @���J  fD9��   tfD9��   ��	  ����E�������	  E1�1��   H�L$pH�AH;A��  H��H�A�����f�D$xH�AH;A�1  � E1�f����  f�|$h�H�L$`��H���� Љ���  A8��z  �S �   H�D$8   ��tHc�H�D$8H��$�   ��HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    �b  ���  D���   ���E���D$X�y  @���	  1��D$^ f�D$\�D$8D�x0H�|$8
A���G  fA��/�l  fE9��b  ��0����V  �T$\�L$Xf9���  �չ��  )�D��A9����A��L$^f�D$\H�L$pH�AH;A��  H��H�A�����f�D$xH�AH;A�  � E1�f����=  f�|$h       �H�L$`��H��A��A ���  A8���  L��$�   A�   M����  E����  @����  H��$0  1�f�H��$(  �    E��tH��$(  �H��$   foT$pH��$�   H�D$@H��H9�t�� H��$   H�ĸ   [^_]A\A]A^A_�f�     ����
��@��D���E��@�ǃ���@��x  H�L$pE1�   H�AH;A�\���H��PPH�L$p�����f�D$xH���P���A�   �c���@ H�L$pD�l$xH��tfA�����  @���S ������     1��X���f�     H�AH;A�B  � 1�f���� ���H�D$`    ������ A�U�f��	�����A�U�f����  ��W���������     L��$�   E1�M���M���L�|$@A��L����r H�SM��H�K��3 ���X  E��u@��tH��$�    ����@�������|$^ �	  H��$0  �����f�H��$(  �    ����f�H�L$p�D$^H�AH;A�K���H��PPH�L$p�����f�D$xH���?���A�   �R���D�l$xH�L$pfA��������H�������H�AH;A��  D�(fA����l���H�D$p    H�|$8
��������  ����@ H�AH;A��  � 1�f��������H�D$`    D�������f�H�AH;A��  D�(fA��������H�D$p    �����D  A���������D  A��AfA���Q�����7�����f�     H�D$p    A�   �����@����  H���   E1��D$^ H�D$HH�D$@fD�|$\H��H�D$P�C ����   fD9kJ��   E��L!      ��$�   ��  H��$�   M�}H;D$P��  H��$�   I9���  F�$(H��$�   E1�L��$�   B�8 H�L$pH�AH;A��   H��A�����H�AfD�T$xH�AH;A��  � E1�f����M  f�|$h�H�L$`��H��A��A ��,  D8���   L��$�   �n���fD  fD;kH����H�D$HH�T$8fD9(tD  H��H�������fD9(u�H+D$H�L$\H���P���O�f9L$X��   H�L$pD�t$^H�AH;A�'���H��PPH�L$pA�����fD�L$xH������E���1���D�l$xH�L$pfA����j���H���a���H�AH;A�-  D�(fA����D���H�D$p    �6�����T$\���  )���D��A9����A��L$^f�D$\�t��� H�AH;A�M  � 1�f��������H�D$`    D������f�H�L$@E1�E1�L��H�D$    �4m H��$�   �����1��������H��$�   HǄ$�       H�D$@H��$�   H��$�   Ƅ$�    H�D$8   f�H�L$@�    �i �����S �D$_ �   1�E1�E1�� �����   �r���fD  H��PH�����D  H��PH����D  H�AH;A��  � 1�f����C���H�D$`    ���3��� H�AH;A��  � 1�f��������H�D$p    ������� H�D$p    A�   �����t$\���؀|$_ D�H��$0  f������H��$(  �    �����     H�AH;A�/  D�(fA��������H�D$p    ����D  �D$_ �&����T$xH��������S A������H�D$p    E������1��"         �����H��PH�����H��PH�����ƿ   ����H��PHA���"���H��PH�N���H��PH����E1�A���D$^ 1�L��$�   fD�D$\�����H��PHA���n���E1�A���D$^ 1�L��$�   fD�\$\����E1�������H��PP����H��PH�m���H��PH�2���H��PHA�������H��PHA�������H��H�D$@H��$�   H��H9�t藀 H����G�����������������AWAVAUATUWVSH���   A�   H��$@  �Ao �Ao	H��$   H���   H��$�   )�$�   )�$�   ����D�vH��A��JA��@tA��A�   �
   DE�f��$�   �H��$�   @��H����@ �����
  f��$�   �H��$�   ��H���� Љ��;
  @8���	  H��$�   D��$�   H��tfA�����
  ���   �S fD9��D$wtfD9��   ��
  ��uifD9cHtrH��$�   H�AH;A��  H��H�AH��$�   �����H��$�   H��f��$�   �O���������
  �S 1�1��  �     fD9cJu�f�     1�1���tfD9cJ�~  fD9cH��  fD9��   �  @���k  fD9��   tfD9��   �W
  A����E������d
  1�1�A�   H��$�   H�AH;A�.  H��A�����H�AfD��$�   H�AH;A��  � E1�f����)  f��$�   �H��$�   ��H���� Љ��  D8���  �S �   H�D$@   A��tIc�H�D$@H��$�   ��HǄ$�       H�D$`H��$�   H��$�   Ƅ$�    ��  H�       ��|$w H���#      �����D���   HE�Ic�H��H�T$P1�H�D$XH��E��H�D$H�{  @���h	  �D$@E1�H�D$8    D�x0H�|$@
A���^  fA��/��  fE9��x  ��0����l  H�T$8H�L$HH9���  H�T$PH�H�L$XH)�H9���HЃ�A	�H�D$8H��$�   H�AH;A�?  H��A�����H�AfD��$�   H�AH;A�j  � E1�f����z  f��$�   �H��$�   ��H��A��A ���  A8��m  L��$�   A�   M����  fD  ����  @����  H��$P  H�     H��$H  �    E��tH��$H  �H��$   fo�$�   H��$�   H�D$`H��H9�t��{ H��$   H���   [^_]A\A]A^A_�fD  ��A��
��@������E��@��A����@��Y  1�A�   ����f�     H��$�   D��$�   H��tfA�����  @���S �f���f�1��F���f�     H��PPH��$�   A�����fD��$�   H�������A�   �����H�AH;A�q  � 1�f��������HǄ$�       �������A�T$�f��	�����A�T$�f����  ��W��������D  L��$�   E1�M���L���L�|$`@��L����e H�SM��H�K��& ����  ��u@��tH��$�    ����@������E���H  H�       ��|$w H��������H��$P  HD�H�H��$H  �    �����A�   ����f�D��$�   H��$�   fA��������H�������H�AH;A��  D� fA����q���H�|$@
HǄ$�       ���$      �����  �����H�AH;A�Y  � 1�f����	���HǄ$�       D�������H�AH;A�?  D� fA��������HǄ$�       ������������� A��AfA���q�����7�����f�     HǄ$�       A�   �����f�     @���  H���   E1�H�D$8    H�D$hH�D$`H��H�D$x�C ����   fD9cJ��   ��L��$�   ��  H��$�   M�|$H;D$x��  H��$�   I9���  B�, H��$�   1�L��$�   B�8 H��$�   H�AH;A�`  H�������H�Af��$�   H�AH;A�  � E1�f�����  f��$�   �H��$�   ��H��A��A ���   D8�utL��$�   �x����    fD;cH����H�D$hH�T$@fD9 tD  H��H�������fD9 u�H+D$hH�L$8H���P���O�H9L$HsbE���!����    H��$�   D��$�   H�������fA��������H�AH;A��  D� fA����m���HǄ$�       �\���H�T$8H�H�T$PH�L$XH)�H9���HЃ�A	�H�D$8����H�AH;A��  � 1�f��������HǄ$�       D�������H�L$`E1�E1�L��H�D$    �r` H��$�   �$���D  H��PPH��$�   A�����fD��$�   H�������A�   �����1�A���_���H��$�   HǄ$�       H�D$`H��$�   H��$�   Ƅ$�    H�D$@   f�     H�L$`�    �\ �I����S �D$w �   1�E1�1������f�H��PPH��$�   �����f��$�   H�������E������@ %      �   �,���fD  H��PH�O���D  H��PH����D  H�AH;A��  � 1�f��������HǄ$�       ������H�AH;A��  � 1�f����T���HǄ$�       ���A���HǄ$�       A�   �o���f�     H�t$8H��H�؀|$w HD�H��$P  H�����H��$H  �    �V���f�     H�AH;A�;  D� fA�������HǄ$�       ����f��D$w ������$�   H�������S A���z���f.�     HǄ$�       E���?���1��   �=���H��PH����H��PH�����ƿ   �*���H��PHA������H��PH�����H��PH����A��E1�1�L��$�   H�D$8    �}���H��PHA������A��L��$�   E1�1�H�D$8    �Q���E1����G���H��PP�W���H��PH�Q���H��PH����H��PHA���>���H��PHA������H��H�D$`H��$�   H��H9�t�Ks H���:�����AWAVAUATUWVSH���   A�   H��$0  �Ao �Ao	H��$  H���   H��$�   )�$�   )L$p謗��D�vH��A��JA��@tA��A�   �
   DE�f��$�   �H��$�   @��H����@ ����2
  f�|$x�H�L$p��H���� Љ���	  @8��_	  H��$�   D��$�   H��tfA����z
  ���   �S fD9��D$otfD9��   ��
  ��ubfD9cHtkH��$�   H�AH;A�O  H��H�AH��$�   �����H�T$pH��f��$�   ���������;
  �S 1�1���   @ fD9cJu�f�     1�1���t&      fD9cJ�.  fD9cH�R  fD9��   ��  @���;  fD9��   tfD9��   �
  A����E������
  1�1�A�   H��$�   H�AH;A��  H��A�����H�AfD��$�   H�AH;A�Y  � E1�f�����  f�|$x�H�L$p��H���� Љ���  A8��b  �S �   H�D$8   A��tIc�H�D$8H��$�   ��HǄ$�       H�D$PH��$�   H��$�   Ƅ$�    �Y  D���   Ic�H������H��H�T$H1�H��H�D$@E���\  @���9	  �D$8E1�H�D$0    D�x0H�|$8
A���N  fA��/�s  fE9��i  ��0����]  H�T$0H�L$@H9���  H�T$HH�H��H��H9���HЃ�A	�H�D$0H��$�   H�AH;A�  H��A�����H�AfD��$�   H�AH;A�=  � E1�f����M  f�|$x�H�L$p��H��A��A ���  A8��V  L��$�   A�   M����  ����  @����  H��$@  H�     H��$8  �    E��tH��$8  �H��$  fo�$�   H��$�   H�D$PH��H9�t��n H��$  H���   [^_]A\A]A^A_�D  ��A��
��@��"���E��@��A����@��F  1�A�   �5���f�     H��$�   D��$�   H��tfA�����  @���S �����f�1��p���f�     H��PPH��$�   A�����fD��$�   H�������A�   ����H�AH;A�Q  � 1�f�������H�D$p    �������f�A�T$�f��	�����A�T$�f����  ��'      W��������fD  L��$�   E1�M���M���L�|$P@��L����X H�SM��H�K�� ���w  ��u@��tH��$�    ����@������E���(  H��$@  H� ����H��$8  �    ����fD  A�   �=���D  D��$�   H��$�   fA��������H�������H�AH;A��  D� fA��������H�|$8
HǄ$�       �������  �����H�AH;A�I  � 1�f���� ���H�D$p    D������H�AH;A�2  D� fA�������HǄ$�       ��������������fD  A��AfA���������7����f�     HǄ$�       A�   � ���f�     @���	  H���   E1�H�D$0    H�D$XH�D$PH��H�D$`�C ����   fD9cJ��   ��L��$�   ��  H��$�   M�|$H;D$`��  H��$�   I9���  B�, H��$�   1�L��$�   B�8 H��$�   H�AH;A�P  H�������H�Af��$�   H�AH;A��  � E1�f�����  f�|$x�H�L$p��H��A��A ���   D8�ujL��$�   ����fD;cH�2���H�D$XH�T$8fD9 tf�H��H������fD9 u�H+D$XH�L$0H���P���O�H9L$@sbE���1����    H��$�   D��$�   H�������fA��������H�AH;A��  D� fA����}���HǄ$�       �l���H�T$0H�H�T$HH��H��H9���HЃ�A	�H�D$0�����H�AH;A��  � 1�f��������H�D$p    D�������f�H�L$PE1�E1�L��H�D$    �(      �S H��$�   �6����    H��PPH��$�   A�����fD��$�   H�������A�   �����1�A�������H��$�   HǄ$�       H�D$PH��$�   H��$�   Ƅ$�    H�D$8   f�     H�L$P�    �O �����S �D$o �   1�E1�1��)���f�H��PPH��$�   �����f��$�   H�������E������@ �   �<���fD  H��PH����D  H��PH����D  H�AH;A��  � 1�f��������H�D$p    ������� H�AH;A��  � 1�f��������HǄ$�       ������HǄ$�       A�   ����f�     H�t$0H��H�؀|$o HD�H��$@  H������H��$8  �    �v���f�     H�AH;A�;  D� fA����i���HǄ$�       �X���f��D$o �������$�   H���ּ���S A�������f.�     HǄ$�       E���O���1��   ����H��PH����H��PH�����ƿ   �t���H��PHA�������H��PH�����H��PH����A��E1�1�L��$�   H�D$0    ����H��PHA������A��L��$�   E1�1�H�D$0    �x���E1����n���H��PP����H��PH�Q���H��PH����H��PHA���>���H��PHA������H��H�D$PH��$�   H��H9�t�kf H����-�����AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`�Պ��D�sH��A��JA��@�P  A��A�
   �@  H�D$pH�T$`H��H�D$(H�T$0��������)      �J  �T$xH�L$(諺�������   f9��F �D$_tf9��   �  ����  f9^H��  H�L$pE1�1��F� �����H�T$0f�L$xH�L$(荹�������6   H�D$8   A��tIc�H�D$8H��$�   1�1�I��H�D$H�@� �~  H��$�   �n  �����1҉�A��D$X���   ���D$^��  E1�@���
  �D$8E1�f�L$@��0f�D$\H�|$8
���;  f��/�a  f9\$\�V  ��0����J  D9t$X��  E���H�L$p��D9���A�A��H�AA	�H;A��  H��H�A�D$@H�T$0H�L$(f�D$x�s���������  H��$�   H�y� ��  fD  E���&  @���  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�� H��$�   H�Ę   [^_]A\A]A^A_��    f9^J����fD  E1�1��t
f9^J�M  f9^H�C  f9��   �  @���-  f9��   tf9��   �D  A����E������;  E1�1�A�   H�L$pH�AH;A�  H�������H�Af�T$xH�AH;A��  � E1�f�����  f�|$h�H�L$`��H���� Љ��  D8���   �   �c��� H�D$pA�   H�T$`H��H�D$(H�T$0辶�����������1�E1�1��D$_ H�D$8   A�   �+���@ ��A��
��@������E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$p�����f�D$xH�������A�   �����    H�L$p�\*      $xH��t
f����W  @����  �F �*���D  H�AH;A�3  � 1�f��������H�D$`    ������ �S�f��	������S�f���F  ��W��������f.�     H��$�   1�H�y� ����L��$�   A��L���w� H�VM��H�N� ����  E��H��$�   u@��tH�y� �����@�������E����  H��$  � ����H��$  �    �����H�L$pA�   H�AH;A�A���H��PP�>���f.�     �T$xH�L$(�q���������f.�     H�AH;A�w  �f��������H�D$p    �����    A��������D  1������f�     ��Af���������7�h���H�D$p    A�   �����    @���  H���   E1�E1�f�L$\H�D$@H��$�   H�D$P�F ��t{f9^JuuE����  H�L$PA����� E1�H�L$pH�AH;A��   H��H�A�D$\H�T$0H�L$(f�D$x藳�������$����T$xH�L$(�>������F ��u�@ f;^H�����H�D$@H�T$8f9t�    H��H�������f9u�H+D$@H���P���O�D9t$Xs%H�L$pD�|$^H�AH;A�T���H��PP�Q����E�����D9���A�A��A	����� A�   ����D  H��$�   �    �� �{���f�     1�E1�1��D$_ �.���H��PH�����@ H��PH�d���D  D���؀|$_ DE�H��$  D�0�A���f�H��$  �    �����T$xH�L$(��������F �s���1��   �����ǽ   ����H��PH����+      ��1ۉ�������E1�1�������E1�E1�1�����H��H��$�   H�T$HH�H���� H���	%�����������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`����D�sH��A��JA��@��  A��A�
   �P  H�D$pH�T$`H��H�D$ H�T$(�4���������  �T$xH�L$ �۱�������   f9��F �D$Xtf9��   �  ����  f9^H�  H�L$pE1�1��v� H�T$(A�����H�L$ fD�L$x軰��������  �H�D$0   A��tIc�H�D$0H��$�   1�1�I��H�D$H�p� �~  H��$�   ��  �D$X1�D�d$\D���   ������D$@A��E���D$8�D$D�K  @����  �D$0A��E1���0f�D$DH�|$0
���p  f��/��  f9\$D��  ��0����  D9t$8�  �T$@E��H�L$p)�D9���A�A��H�AA	�H;A�   H��H�AH�T$(�����H�L$ f�D$x薯��������  H��$�   H�y� �  f�     E���V  @���L  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�#� H��$�   H�Ę   [^_]A\A]A^A_��    f9^J�����fD  E1�1��t
f9^J�}  f9^H�s  f9��   �6  @���]  f9��   tf9��   ��  A����E�������  E1�1�A�   H�L$pH�AH;A�4  H��A�����H�AfD�D$xH�AH;A�  � E1�f����  f�|$h�H�L$`��H���� Љ��,      D  A8��  �   �Q����H�D$pA�   H�T$`H��H�D$ H�T$(�ޭ�����������H��$�   1�1�I��H�D$H�� �~ H��$�   @���  D���   1��D$X E��D���t  E1�E1��������A��
��@������E��@��A����@���  H�L$pE1�A�   H�AH;A�����f.�     H��PPH�L$p�����f�T$xH�������A�   ������    H�L$p�\$xH��t
f����W  @����  �F �����D  H�AH;A�s  � 1�f��������H�D$`    ������ �S�f��	������S�f���F  ��W��������f.�     H��$�   1�H�y� �����L��$�   A��L���g� H�VM��H�N� ���  E��H��$�   u@��tH�y� �����@�������E����  �D$XH��$  ������H��$  �    ����fD  H�L$pA�   H�AH;A� ���H��PP������T$xH�L$ �]������w���fD  H�AH;A��  �f��������H�D$p    �����    A���������D  1�����f�     ��Af���������7�3���H�D$p    A�   �����E1�1�H�D$0   �D$D����D$@����D$\   �@���2  H���   E1�E1�H�D$8H��$�   A�����H�D$P�F ��tzf9^JutE����  H�L$PA���� E1�H�L$pH�AH;A��   H��H�AH�T$(fD�d$xH�L$ �j�������������T$xH�L$ �������F ��u��    f;^H�����H�D$8H�T$0f9t�    -      H��H�������f9u�H+D$8H���P���O�D;t$Dv%H�L$pA�   H�AH;A�U���H��PP�R�����T$@D�t$\)�D9���A�A��A	�����A�   �T���1�E1�1��D$X H�D$0   A�   f�     H��$�   �    �>� �����f�     1�E1�1��D$X ����H��PH����@ H��PH�����D  D���؀|$X DE�H��$  D�0�����f�H��$  �    ������T$xH�L$ 让�����F ����1��   �'����ǽ   �*���H��PH���?���1ۉ��)�����E1�E1�1�������E1�1�����H��H��$�   H�T$HH�H��� H��������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`�x��D�sH��A��JA��@�P  A��A�
   �@  H�D$pH�T$`H��H�D$(H�T$0���������J  �T$xH�L$(苨�������   f9��F �D$_tf9��   �  ����  f9^H��  H�L$pE1�1��&� �����H�T$0f�L$xH�L$(�m��������6   H�D$8   A��tIc�H�D$8H��$�   1�1�I��H�D$H� � �~  H��$�   �n  �����1҉�A��D$X���   ���D$^��  E1�@���
  �D$8E1�f�L$@��0f�D$\H�|$8
���;  f��/�a  f9\$\�V  ��0����J  D9t$X��  E���H�L$p��D9���A�A��H�AA	�H;A��  H��H�A�D$@H�T$0H�L$(f�D$x�S���������  H��$�   H�y� ��  fD  E���& .       @���  H��$  �     H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p��� H��$�   H�Ę   [^_]A\A]A^A_��    f9^J����fD  E1�1��t
f9^J�M  f9^H�C  f9��   �  @���-  f9��   tf9��   �D  A����E������;  E1�1�A�   H�L$pH�AH;A�  H�������H�Af�T$xH�AH;A��  � E1�f�����  f�|$h�H�L$`��H���� Љ��  D8���   �   �c��� H�D$pA�   H�T$`H��H�D$(H�T$0螤�����������1�E1�1��D$_ H�D$8   A�   �+���@ ��A��
��@������E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$p�����f�D$xH�������A�   �����    H�L$p�\$xH��t
f����W  @����  �F �*���D  H�AH;A�3  � 1�f��������H�D$`    ������ �S�f��	������S�f���F  ��W��������f.�     H��$�   1�H�y� ����L��$�   A��L���W� H�VM��H�N�� ����  E��H��$�   u@��tH�y� �����@�������E����  H��$  � ����H��$  �    �����H�L$pA�   H�AH;A�A���H��PP�>���f.�     �T$xH�L$(�Q���������f.�     H�AH;A�w  �f��������H�D$p    �����    A��������D  1������f�     /      ��Af���������7�h���H�D$p    A�   �����    @���  H���   E1�E1�f�L$\H�D$@H��$�   H�D$P�F ��t{f9^JuuE����  H�L$PA����� E1�H�L$pH�AH;A��   H��H�A�D$\H�T$0H�L$(f�D$x�w��������$����T$xH�L$(�������F ��u�@ f;^H�����H�D$@H�T$8f9t�    H��H�������f9u�H+D$@H���P���O�D9t$Xs%H�L$pD�|$^H�AH;A�T���H��PP�Q����E�����D9���A�A��A	����� A�   ����D  H��$�   �    �n� �{���f�     1�E1�1��D$_ �.���H��PH�����@ H��PH�d���D  D���؀|$_ DE�H��$  D�0�A���f�H��$  �    �����T$xH�L$(�ޠ�����F �s���1��   �����ǽ   ����H��PH������1ۉ�������E1�1�������E1�E1�1�����H��H��$�   H�T$HH�H���� H���������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H��$�   H���   H��$�   )D$p)L$`��o��D�sH��A��JA��@�S  A��A�
   �@  H�D$pH�T$`H��H�D$(H�T$0���������J  �T$xH�L$(軟�������   f9��F �D$_tf9��   �  ����  f9^H��  H�L$p�����E1��S| H�T$0f�l$x1�H�L$(蝞�������6   H�D$8   A��tIc�H�D$8H��$�   1�1�I��H�D$H�P� �~  H��$�   �n  ���  �A���D$X���   ��0      �D$^��  E1�@���  �D$8E1���0f�D$@H�|$8
���C  f��/�i  f9\$@�^  ��0����R  fD9t$X��  E�����  )�A��9�H�L$p��A�A��A	�H�AH;A��  H��H�AH�T$0A�����H�L$(fD�T$x肝��������  H��$�   H�y� ��  D  E���&  @���  H��$  E1�fD� H��$  �    ��tH��$  �H��$�   H��H�T$HfoT$p�� H��$�   H�Ę   [^_]A\A]A^A_�fD  f9^J����fD  E1�1��t
f9^J�M  f9^H�C  f9��   �  @���-  f9��   tf9��   �D  A����E������;  E1�1�A�   H�L$pH�AH;A�  H�������H�Af�|$xH�AH;A��  � E1�f�����  f�|$h�H�L$`��H���� Љ��  D8���   �   �c��� H�D$pA�   H�T$`H��H�D$(H�T$0�Λ�����������1�E1�1��D$_ H�D$8   A�   �+���@ ��A��
��@������E��@��A����@���  H�L$pE1�A�   H�AH;A����f.�     H��PPH�L$pA�����fD�\$xH�������A�   ����D  H�L$p�\$xH��t
f����W  @����  �F �*���D  H�AH;A�3  � 1�f��������H�D$`    ������ �S�f��	������S�f���F  ��W��������f.�     H��$�   1�H�y� ����L��$�   A��L���� H�VM��H�N�� ����  E��H��$�   u@�1      �tH�y� �����@�������E����  H��$  �����f�H��$  �    �����H�L$pA�   H�AH;A�>���H��PP�;����     �T$xH�L$(聚��������f.�     H�AH;A�w  �f��������H�D$p    �����    A��������D  1������f�     ��Af���������7�`���H�D$p    A�   �����    @���  H���   E1�E1�H�D$@H��$�   H�D$P�F ���|   f9^JuvE����  H�L$PA����� E1�H�L$pH�AH;A��   H��H�AH�T$0A�����H�L$(fD�L$x覘�������$����T$xH�L$(�M������F ��u� f;^H�����H�D$@H�T$8f9t�    H��H�������f9u�H+D$@H���P���O�fD9t$Xs$H�L$pD�|$^H�AH;A�R���H��PP�O���E�����  )�A��9���A�A��A	�����A�   ����f�H��$�   �    �� �{���f�     1�E1�1��D$_ �.���H��PH�����@ H��PH�d���D  D���؀|$_ DE�H��$  fD�0�A����H��$  �    �����T$xH�L$(�������F �s���1��   �����ǽ   ����H��PH������1ۉ�������E1�1�������E1�E1�1�����H��H��$�   H�T$HH�H��� H���
�����������AWAVAUATUWVSH��   H��$  �Ao �Ao	H��$�   H���   H��$�   )�$�   )L$p�g��D�kH��A��JA��@��  A��A�
   ��  H��$�   H�T$pH��H�D$ 2      H�T$(�>��������  ��$�   H�L$ ���������   f9��F �D$_tf9��   �>  ���&  f9^H�,  H��$�   E1�1��zs H�T$(A�����fD��$�   H�L$ 輕��������  f�H�D$0   A��tIc�H�D$0H��$�   1�1�I��H�D$`�p� �~  H��$�   �  H�       ��|$_ H��������HE�Ic�D���   H��H�T$81�H�D$@H��I��H�D$PE���d  @����  �D$0A��E1��0f�D$HH�|$0
���x  f��/��  f9\$H��  ��0�����  M9��.  L�l$8H�H�T$@H)�L9���I�A��A	�H��$�   H�AH;A�  H��H�AH�T$(�����H�L$ f��$�   �t���������  H��$�   H�y� �  �    E���V  @���L  H��$   H�     H��$  �    ��tH��$  �H��$�   H��H�T$`fo�$�   ��� H��$�   H�Ĩ   [^_]A\A]A^A_� f9^J�����fD  E1�1��t
f9^J�}  f9^H�s  f9��   �F  @���]  f9��   tf9��   ��  A����E�������  E1�1�A�   H��$�   H�AH;A�b  H��A�����H�AfD��$�   H�AH;A�  � E1�f����  f�|$x�H�L$p��H���� Љ��>  A8���   �   �+���H��$�   A�   H�T$pH��H�D$ H�T$(趒�������x���H��$�   1�1�I��H�D$`胲 �~ H��$�   @���	  D���   1��D$_ E��D���o  E1�E1�������     3      ��A��
��@������E��@��A����@���  E1�A�   ������     H��$�   ��$�   H��t
f�����  @����  �F �$���H��PPH��$�   �����f��$�   H�������A�   ����H�AH;A��  � 1�f��������H�D$p    ������ �S�f��	������S�f���F  ��W��������f.�     H��$�   1�H�y� �����L��$�   A��L���G� H�VM��H�N�w� ���?  E��H��$�   u@��tH�y� �����@�������E����  H�       ��|$_ H��������H��$   HD�H�H��$  �    ����@ A�   �����D  ��$�   H�L$ �>������p����    H�AH;A��  �f����d���HǄ$�       �S���@ A���������D  1��y���f�     ��Af���������7�+���HǄ$�       A�   �����H��������E1�1�H�D$0   H�D$PH��������H�D$@H�D$8   @���D  H���   E1�E1�H�D$HH��$�   A�����H�D$h�F ��t|f9^JuvE����  H�L$hA���� E1�H��$�   H�AH;A�#  H��H�AfD��$�   H�T$(H�L$ �3��������������$�   H�L$ �׏�����F ��u�f;^H�����H�D$HH�T$0f9t@ H��H�������f9u�H+D$HH���P���O�L;l$PvA�   �Q���f.�     L�l$8H�H�T$@H)�L9���I�A��A	��"���H��PP�����A�   ����1�E1�1��D$_ H�D$0   A�   f.4      �     H��$�   �    �� �����f�     H��PP�����D  1�E1�1��D$_ �n���H��PH�e���@ H��PH�����D  L��H�؀|$_ LE�H��$   L�(�����H��$  �    ������$�   H�L$ �k������F �����1��   ������ǽ   �����H��PH������1ۉ�������E1�E1�1��������E1�1������H��H��$�   H�T$`H�H��N� H���v ��������AWAVAUATUWVSH��   H��$  �Ao �Ao	H��$�   H���   H��$�   )�$�   )L$p�r]��D�sH��A��JA��@�M  A��A�
   �`  H��$�   H�T$pH��H�D$(H�T$0螌�������T  ��$�   H�L$(�B��������   f9��F �D$otf9��   �  ���  f9^H�  H��$�   E1�1���i �����H�T$0f��$�   H�L$(���������7  @ H�D$8   A��tIc�H�D$8H��$�   1�1�I��H�D$X�Ы �~  H��$�   �^  D���   Ic�H������1�I��H�D$HH��I��H�D$@E����  E1�@���   �D$8E1�A�σ�0f�D$PH�|$8
���0  f��/�V  f9\$P�K  ��0����?  L9l$@��  L�l$HH�H��H��L9���I�A��A	�H��$�   H�AH;A��  H��H�AfD��$�   H�T$0H�L$(����������v  H��$�   H�y� ��   E���  @���  H��$   H�     H��$  �    ��tH��$  �H��$�   H��H�T$Xfo�$�   �� H��$�   H�Ĩ   5      [^_]A\A]A^A_� f9^J�����fD  E1�1��t
f9^J�  f9^H�  f9��   �  @����  f9��   tf9��   �7  A����E������.  E1�1�A�   H��$�   H�AH;A�"  H�������H�Af��$�   H�AH;A�~  � E1�f�����  f�|$x�H�L$p��H���� Љ��   D8���   �   �M���H��$�   A�   H�T$pH��H�D$(H�T$0�8������������1�E1�1��D$o H�D$8   A�   ������A��
��@������E��@��A����@���  E1�A�   �����fD  H��$�   ��$�   H��t
f����a  @����  �F �d���H��PPH��$�   �����f��$�   H�������A�   �����H�AH;A�3  � 1�f��������H�D$p    ������� �S�f��	������S�f���&  ��W��������f.�     H��$�   1�H�y� �+���L��$�   A��L���� H�VM��H�N�7� ����  E��H��$�   u@��tH�y� �����@�������E����  H��$   H� ����H��$  �    �����A�   �L���f���$�   H�L$(������������    H�AH;A��  �f��������HǄ$�       �s���@ A�����>���D  1������f�     ��Af���������7����HǄ$�       A�   �F���@ @���A  H���   E1�E1�f�L$lH�D$PH��$�   H�D$`�F ����   f9^J�~   E����  H�L$`A��薽 E1�H��$�   H�A6      H;A�  H��H�A�D$lH�T$0H�L$(f��$�   �9��������I�����$�   H�L$(�݆�����F ���x���f;^H�����H�D$PH�T$8f9tfD  H��H�������f9u�H+D$PH���P���O�L9l$@sE���J���L�l$HH�H��H��L9���I�A��A	��'���f.�     H��PP�}���D  A�   ����D  H��$�   �    �.� ����f�     H��PP�����D  1�E1�1��D$o �.���H��PH�����@ H��PH�z���D  L��H�؀|$o LE�H��$   L�(�Q����H��$  �    ������$�   H�L$(苅�����F ����1��   �����ǽ   ����H��PH���\���1ۉ�������E1�1�������E1�E1�1�����H��H��$�   H�T$XH�H��n� H������������AWAVAUATUWVSH��   H��$�   �Ao �Ao	H��$�   H���   H�L$v)D$`)L$PH�l$`�T��H��H��H�D$PH��H�D$(�������(  ��1�E1�E1�f�     H�D$w1�1�I��H�D$H誣 �~  H�D$x��  ���   ���D$7�H  @���b  E1�A������C���f��	wz��0���trH��$   ��0���� A�   H�L$`H�AH;A�^  H��H�AH�T$(H��fD�|$h�+�������  �T$hH���փ���ÍC���f��	v��     f9^H��  f9��   tf9��   �N  D����A ��?  H��$   �e   �߹ H�L$`H�AH;A��  H��H�AH�T$(H��fD�|$h葂������  �T$hH���<���f9��   ���]7        f9��   �-   �P  E������� @���  H���   E1�H�D$8�F H�T$xL���   H�T$@ ��t
f9^J��  f9^H�  H�\$xA�H�C���  H��tH�L$@A���� H��$   �.   �� �|$7H�L$`H�AH;A�  H��H�AH�T$(�����H��f�D$h蚁�����b  H�\$xH�C�H��tB@��uxE��usL�t$xA��L��艸 H�\$xH�VM��H�N�� ��uH��$�   �    H��$�   H�K�H�T$HfoT$`�3� H��$�   H�Ĉ   [^_]A\A]A^A_�L�t$x�H�D$8f9�  H��L9�u�f9��   tf9��   �A���H�\$xD���A �H�C��2���H��t	@����  H��$   �e   軷 H�L$`�1^ �����H��f�T$hH�T$(�z������v  �T$hH���%������   ���F f9��  f9��   �  E������f.�     �T$hH���������F ������     �+   H��$   �� H�L$`E��H�AH;A�����H��PP����H+D$8H��$   H���P0���� H�L$`A��D�d$7H�AH;A�����H��PP�����f.�     D��o  E���0  H�L$@A��萶 E1�E1�����D  ��D��_���H��$   �.   �c� E1��   �����fD  ��t
f9^J�@  f9^H�����f9�H��$   ���ҍT+�� E���*���fD  H�L$@A���� �0���H��PP�.���L�t$x�    L��萳 �����T$hH���n�����   ���F f9���   f9��   ��   E1�E1�A�������t
f9^8      J��   f9^H��   f9��   ��   E��tEH�L$`A��H�AH;AsdH��H�AH�T$(H��fD�t$h�'~����t'��A���I���f�     H��$   �0   �� ��T$hH��A�   �~�����F �_���H��PP�fD  1��������t
f9^J�0���f9^H�&���f9�H��$   ��E1�E1��ҍT+豴 H�L$`�'[ H�T$(�����f�L$hH���p}������������T$hH���~�����F �����H��$   E1�1�H��$   H� L�@��� H�\$xH�{� ����������H�\$xH�C�L�t$xH�����������H�\$xL�t$xH�{� ���������A��A������H��H�D$xH�T$HH�H��Ѡ H����������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P`H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PPH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PXH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PHH��H��`[ÐSH��`L�$  H��Ao�Ao	L��$�   H�@(H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H9      �L$ H��L�L$0L�L$@u�ؿ��H��H��`[���H��H��`[Ð���SH��`L�  H��Ao�Ao	L��$�   H�@H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u�(���H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@0H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u�����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@ H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u�H���H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@8H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���SH��`L��  H��Ao�Ao	L��$�   H�@@H��)\$PH��$�   )L$@L��$�   L�D$(L�D$PL9�H�L$ H��L�L$0L�L$@u����H��H��`[���H��H��`[Ð���WVSH��   H��$�   �Ao�Ao�{)T$PL�L$PH��H��$�   )L$@L�D$`���ᵃ��KH�L$pH�D$0H��$�   H�\$ )L$`H�D$(�1���H�D$pH��$�   H�D$@H��$�   foD$@f�D$x�{H�H��H�Đ   [^_Ð��AWAVAUATUWVSH��   H��$   M�QM�(M�pM�	H���@L��$�   L��$�   L��$�   L��$�   ��   H��$(  L�L$PH�L$pL��$�   H�D$ L�D$0L�L$PL�D$`L�l$`H�\$(Ǆ$�   ���:      �L�t$hL�T$X����H�D$pH��$�   �D$xf��$�   ��$�   ����  H��$0  ��#fo�$�   H��H�ĸ   [^_]A\A]A^A_�H���   A�   A�   H��$�   A������F��H�x@ I��A��H�x0 @��1ېA���  f��$�   �H��$�   @��H����@ �����  f��$�   �H��$�   ��H���� �A���}  @8���  ��$�   H��$�   f���u	H����  H�E����   I�W8�Zf9�A���%  @���9  I�W(f9
A��D��D��Q  H��$�   H��H�AH;A��  H��H�AfD��$�   E����   I9_@A��E����   D��A�������1�E��tI9_@u	H���|  E��tI9_0u	H����  H��$0  ��� ��  H��$(  �    �?���I�W(�Zf9�A���>���E����  I9_@�g  H���^  H��$0  �  1�f�H��$(  �������A��I9_0A��@���=���@������������H�AH;A�q  � 1�f����f���HǄ$�       D��@8��W���f.�     �   �����fD  H�AH;A�  � 1�f��������HǄ$�       �������H�AH;A�  � f�������HǄ$�       � ���@ H��$0  H��$�   H��$�   � H��$(  �    �2s���������H��$(  ������f.�     H��PP����D  E��t+I9_0��   H��$0  �  H��$(  �    ���� H��$0  �  H��$(  �    �q���f�H�D�L$O�T$N�PHD�L$O�T$N������;      H�D�\$OD�L$N�PHD�\$OD�L$N�q���H�D�L$N�PHD�L$N�����H���_���H��$0  � 1������H��$0  E��� t
I9_0�>�����������H��$0  ��鐐�����������AWAVAUATUWVSH��   �AoM�)M�qH��$  H��$�   I��H��)L$@1�1�I��誑 H��$�   �    H��H��$�   �m� H��$  H��$�   H�\$0H��foT$@H�t$(L�L$`L�D$pL�l$`)T$pH�D$ L�t$h����H��$�   H�D$@foD$@fĄ$�   )D$Pfo\$PH�|$P)\$@�\$X�+� H��$   I��I��H��$�   H��$�   �X� f�����H���� �A����   fA�����M���t��uM8�u�H��$�   H�|$@�����fod$@A$$��A���~@L��H�Ĩ   [^_]A\A]A^A_�f�     I�EI;EsV� f������f.�     H��H���T� �f�H�GH;Gs6� f����    �    AD�HD��H����     I�E L���PH�@ H�H���PH��H��H��$�   H��H�H���� H���&���������AWAVAUATUWVSH��   �AoM�)M�qH��$  H��$�   I��H��)L$@1�1�I��芏 H��$�   �    H��H��$�   �M� H��$  H��$�   H�\$0H��foT$@H�t$(L�L$`L�D$pL�l$`)T$pH�D$ L�t$h�����H��$�   H�D$@foD$@fĄ$�   )D$Pfo\$PH�|$P)\$@�\$X�� H��$   I��I��H��$�   H��$�   �H� f�����H���� �A����   fA�����M���t��uM8�u�H��$�   H�|$@�<      ����fod$@A$$��A���~@L��H�Ĩ   [^_]A\A]A^A_�f�     I�EI;EsV� f������f.�     H��H���4� �f�H�GH;Gs6� f����    �    AD�HD��H����     I�E L���PH�@ H�H���PH��H��H��$�   H��H�H��ޑ H������������AWAVAUATUWVSH��   �AoM�)M�qH��$  H��$�   I��H��)L$@1�1�I���j� H��$�   �    H��H��$�   �-� H��$  H��$�   H�\$0H��foT$@H�t$(L�L$`L�D$pL�l$`)T$pH�D$ L�t$h�����H��$�   H�D$@foD$@fĄ$�   )D$Pfo\$PH�|$P)\$@�\$X��� H��$   I��I��H��$�   H��$�   �H� f�����H���� �A����   fA�����M���t��uM8�u�H��$�   H�|$@�����fod$@A$$��A���~@L��H�Ĩ   [^_]A\A]A^A_�f�     I�EI;EsV� f������f.�     H��H���� �f�H�GH;Gs6� f����    �    AD�HD��H����     I�E L���PH�@ H�H���PH��H��H��$�   H��H�H�辏 H�������������SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ 辰��H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �.���H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(=      H��$�   H�D$ ����H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ ����H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �����H��H��`[Ð����SH��`H��$�   �Ao�AoH�D$0H��$�   H��L�L$@)D$@L�D$P)L$PH�D$(H��$�   H�D$ �>���H��H��`[Ð����VSH��8H��$�   H��$�   H�t$xHcI��A��M��H�L$ M��H�H��H�D$(�p� H)��H��8[^Ð���UAWAVAUATWVSH��XH��$�   �E@M�0M�xI���   L��I�͉E�H�M��e8���wH�� L�@JI�ċUHL�\$0����J��@�E��Ã���!Å��ڄ�DUH��A��L�]��D$ I�K薭 L�]�A�   Hc�A)�Mc�M�A�|$  ��   ���7  �UH����   ��   uYH�wHc�H9�|iE��H�G    D��uI�I��L��L���P`H9ظ   E�L��M�u A�uH�e�[^_A\A]A^A_]��    A�D$K��I��H�wHc�A�H9�}�H�FH��������U�H)�H��L�d$0H�\$(Hc�H�t$ M���ӟ M���^���A�D$J��I��A��=���fD  �AH�H�D H�������M�D$A�T$IH)�I�D$L�L�\$2H�L$(L�L$ L��L�]�I��良 L�]���D)ل�M���������   ������EH��������}�@t/����I��A��A��A�BH�A�DJA�AA�D$NA�����A�D$N��I��A��{�������UAWAVAUATWVSH��XH��$�   >      �E@M�(M�xI���   L��I�̉E�H�M��6��D�sH�� �UHL�\$0H��H�L$DL�]�L�GJD��E���J��@�E�@�ƃ���!�@�ƉD$ �M� L�]�A�   Hc�A)�Mc�Mـ  ua@����   H�{Hc�H9���   E��H�C    D��uI�E I��L��L���P`H9Ƹ   E�L��M�,$A�\$H�e�[^_A\A]A^A_]ÍAH�H�D H��������L�G�WIH)�H�GL�L�\$2H�L$(L�L$ L��L�]�I���ͭ L�]���D)�@��M���P���A��   �C����EH���8����}�@tcA����I��A��A�FH��DJA�A�GNA�����H�GH����c����U�H)�H��L�t$0H�t$(Hc�H�|$ M���� M��������GN��I��A���������UAWAVAUATWVSH��XH��$�   �E@M�0M�xI���   L��I�͉E�H�M��%4���wH��0L�@JI��H�UHL�\$0����J��@�E��Ã���!�H��
H�ڄ�HDUH��A��L�]��D$ I�K(�� L�]�A�(   Hc�A)�Mc�M�A�|$  ��   ���3  H�}H ��   ��   uUH�wHc�H9�|eE��H�G    D��uI�I��L��L���P`H9ظ   E�L��M�u A�uH�e�[^_A\A]A^A_]� A�D$K��I��H�wHc�A�H9�}�H�FH���������U�H)�H��L�d$0H�\$(Hc�H�t$ M��蓛 M���b���A�D$J��I��A��A���fD  �AH�H�D H����}���M�D$A�T$IH)�I�D$L�L�\$2H�L$(L�L$ L��L�]�I���I� L�]���D)ل�M���������   �����H�}H ������}�@t/����I��A��A��A�BH�A?      �DJA�AA�D$NA�����A�D$N��I��A���������UAWAVAUATWVSH��XH��$�   �E@M�(M�xI���   L��I�̉E�H�M���1��D�sH��0H�UHL�\$0H��H�L$XL�]�L�GJD��E���J��@�E�@�ƃ���!�@�ƉD$ �̧ L�]�A�(   Hc�A)�Mc�Mـ  ua@����   H�{Hc�H9���   E��H�C    D��uI�E I��L��L���P`H9Ƹ   E�L��M�,$A�\$H�e�[^_A\A]A^A_]ÍAH�H�D H�������L�G�WIH)�H�GL�L�\$2H�L$(L�L$ L��L�]�I��茩 L�]���D)�@��M���P���A��   �C���H�}H �8����}�@tcA����I��A��A�FH��DJA�A�GNA�����H�GH����"����U�H)�H��L�t$0H�t$(Hc�H�|$ M���ޘ M��������GN��I��A��������UWVSH��8H��$�   H��$�   H��$�   H��$�   H��I��A��t]H��M��H�D$ M��H)�Hc�H�H�L$(H��舨 D�1�H��H)�H��A)�Mc�M��u�:�H��8[^_]ÐH��H���E{���)���HcM��H�D$ M��H�H�L$(H���1� )��H��8[^_]Ð���UAWAVAUATWVSH��   H��$�   )u ���   ���   M�(M�p�E�I���   L�����   H�M`H�M�H�UhL�}�H��H�E���.��H�{D��L��I��H�ٸ   H��HH���� �CH��0H�t$@%  =  ��  �:� H�|$ M��H��H�E�H�E�A�-   �t$(H��H�E��߭ ��,�E��  H�M��� LcU�I��I�BH����&���H)�A�C8H�|$@I��<�  ����@        I�H��p��H�@8H9���  M��H��H����y��LcU�M��M����   M�к.   H��D�M�L�U��y��L�U�H��D�M��H  H)�H�A�D$H�A�|$  ��   H�{L��I9��B  E��H�C    D��uI�E I��L��L���P`H9�   E�H�E`L�(�X(u H�e[^_A\A]A^A_]� D�@Ic�D�E�H��H�������H)���� D�E�H�t$@�t$(H�M�H�|$ M��H��H�E��y� �E������A�|$  �G���1�K�DH�����������+H)�H�D$@���   ��  �A�q��u�L��   L�X�E�L$IL�U�H�E�M�D$I�T$H�L$ H�MhL�T$8L�|$0L�\$(�|���u�H�{H�E�Lc�I9�D�U�L��I�������H�GH����.����U�H)�M��H��L�d$@L�T$(Hc�H�|$ M��M���� �}������� H�}�M��H���t$ A�-   H��H�E��e� ��,�E������D�@Ic�D�E�H��H�������H)��i� D�E�M��H��H�t$@�t$ H��H�E��� �E��=���L��L�U�L�]��l��L�U�L�]��]��� A�|$  �����A���v����F<9������N�QЀ�	�����</�����1��M���I��1�����D  I��H��L��N���LcU�M������D  M��H��H��D�U�L�U���v��L�U�D�M�������������������UAWAVAUATWVSH��   H��$�   ���   ���   M�(M�p�E�H���   L�}L��H�MpH�MH�Ux�(I���   H��H�E��}��*��H�{D��L��I��H�ٸ   H��HH�蛚 �CH��@H�t$@%  =  ��  �ڿ H�MM��H��A      �m�H�EA�6   H�|$ H�E�H�M�H�D$(�}�H�E��u� ��5�E�  H�M�� � LcUI��I�BH�������H)�A�C8H�|$@I��<�4  ����  I�H�Rl��H�@8H9���  M��H��H���gu��LcUM��M����   M�к.   H��D�M�L�U��Ou��L�U�H��D�M��^  H)�H�A�D$H�A�|$  ��   H�{L��I9��H  E��H�C    D��uI�E I��L��L���P`H9�   E�H�EpL�(�XH�e([^_A\A]A^A_]�D�@Ic�D�E�H��H�������H)��m� D�E�H�t$@M��H�EH�E�H��H�M�H�|$ �m�H�D$(�}��� �E����D  A�|$  �A���1�K�DH����T������+H)�H�D$@���   ��  �A�q��uL��   L�X�E�L$IL�UH�E�M�D$I�T$H�L$ H�MxL�T$8L�|$0L�\$(����uH�{H�E�Lc�I9�D�UL��I�������H�GH��������U�H)�M��H��L�d$@L�T$(Hc�H�|$ M��M���t� �}�y����G� H�}�M��H���m�H�EA�6   H�|$ H�EH��H�E��}��� ��5�E�s���D�@Ic�D�E�H��H����4���H)��� D�E�H�t$@M��H�M�H�|$ H���m�H�E�}�蕦 �E�$���L��L�U�L�]��g��L�U�L�]��D���A�|$  �����A���f����F<9������V��0��	�����</�����1��=���I��1��t���D  I��H��L��N���LcUM������D  M��H��H��D�U�L�U��Jr��L�U�D�M�������������������SH��@�Ao H�)D$0L�D$0H��H�L$xH�L$(�L$B      p�L$ H���PHH��H��@[Ð���SH��@�Ao H�)D$0L�D$0H���L$x�L$(�L$p�L$ H���PH��H��@[Ð����SH��@H��Ao�D$x)L$0L�D$0H���L$p�D$(�L$ H���P8H��H��@[Ð�SH��PH��$�   �Ao �(H��)D$@H�L$0H�H�L$(��$�   L�D$@�|$0�L$ H���P@H��H��P[Ð��SH��@L��  H��AoD�D$xH�@H��)L$0�L$pD�D$(L�D$0L9ЉL$ H��u����H��H��@[�f���H��H��@[Ð����SH��@L��  H��AoD�D$xH�@ H��)L$0�L$pD�D$(L�D$0L9ЉL$ H��u�{���H��H��@[�f���H��H��@[Ð����SH��@L��  H��AoL�D$xH�@(H��)L$0�L$pL�D$(L�D$0L9ЉL$ H��u����H��H��@[�f���H��H��@[Ð����SH��@L�d  H��AoL�D$xH�@0H��)L$0�L$pL�D$(L�D$0L9ЉL$ H��u�����H��H��@[�f���H��H��@[Ð����VSH��8H��$�   HcL��L��L�D$ L�L$x��L�D$pH�D$(�]� �3H��8[^Ð���UWVSH��XI� I�XA�iH�D$0L�D$0H��L��H��$�   H�\$80ۉ�ᵿ����  H�D$(��$�   A�IH�L$@�D$ �A���H�D$@�n�T$HH�H��H	�H�_H��X[^_]Ð�������������UAWAVAUATWVSH��   H��$�   E�qI�0I�XD���   A��H��M��D���   uPE��E��H��H�u�D�D$ L�E�D�l$(H�]������]H�u �؈�H��H�7H�_H�e([^_A\A]A^A_]�@ I���   D�E�A��H�M�y"��E��D�E�t@Lch0M�L$L�X(M9�C      |@I�D$    E��uH�M��L��H���P`I9�A��D����� Lch@M�L$L�X8M9�}�M)�L�]�I�AH��������H)�A��M��L�M�H�L$0A��   H�M��m��A�� L�M�I�D$    L�]�t4E��L�]�Mc�u�H�M��H��H�U��P`L�]�I9��W���A�   �b���E���Y���H�M��L��H���P`L�M�I9�u�H�Mc�H��M��H�U��P`L9�A���"���������������SH��P��$�   ��$�   �Ao�D$ L�D$@H���D$0�D$(    )L$@����H��H��P[Ð�������SH��`H��$�   �Ao �(H��)D$P�D$(L   H�D$@H�D$0��$�   L�D$P�|$@�D$ ����H��H��`[Ð��������������SH��@�D$x�Ao �D$(�D$pH��L�D$0)D$0�D$ �����H��H��@[Ð���������SH��@�D$x�Ao �D$(�D$pH��L�D$0)D$0�D$ �����H��H��@[Ð���������SH��@H�D$x�Ao H�D$(�D$pH��L�D$0)D$0�D$ ����H��H��@[Ð�������SH��@H�D$x�Ao H�D$(�D$pH��L�D$0)D$0�D$ ����H��H��@[Ð�������VSH��8H��$�   H��$�   H�t$xH��A��LcH�D$ N�HL�L$(M��I��H��蟙 H)�H���H��8[^�UAWAVAUATWVSH��XH��$�   �E@M�0M�xI���   L��I�͉E�H�M�� ���wH��0�UHL�\$0I�ĉ���J��@�E��Ã���!Å��ڄ�DUH��A��L�]��D$ I�K(M�D$L�ŕ L�]�Hcȸ   )�A�|$  H�M�C��   ���P  �UH����   ��   uZH�wHc�H9�|kE��H�G    D��uI�I��D      L��L���P`H9ظ   E�L��M�u A�uH�e�[^_A\A]A^A_]��     A�D$N��I��H�wHc�fA�H9�}�H�D6H����Ž���U�H)�H��L�d$0H�\$(Hc�H�t$ M���1� M���[���f�     A�D$L��I��fA��0���f.�     �AH�H��   H����Z���M�D$A�T$JI�IH)�I�D$L�\$4H�L$(L�L$ L��L�]�I��襗 L�]�L)�M��H��H�����������   ������EH��������}�@t4����I��A��I�t$LA��A�BH��FfA�AA�D$TfA��r���A�D$T��I��fA��\���������UAWAVAUATWVSH��hH��$�   �EPM�(M�xI���   L��I�̉E�H�M����D�sH��0L�@LH�ǋUXL�\$0L�E�H�L$XL�]�D��E���J��@�E�@�ƃ���!�@�ƉD$ �Y� �   L�]�Hc�)ʀ  Hc�M�Sua@����   H�{Hc�H9���   E��H�C    D��uI�E I��L��L���P`H9Ƹ   E�L��M�,$A�\$H�e�[^_A\A]A^A_]ÍAH�H��   H���臻��L�G�WJI�IH)�H�GL�\$4H�L$(L�L$ L��L�]�I���֕ L�]�L)�M��H��H��@���H���A��   �;����EX���0����}�@tiA��H�u���I��A��A�FH��FfA�A�GTfA������H�D?H��������U�H)�H��L�t$0H�t$(Hc�H�|$ M���N� M��������GT��I��fA�������UAWAVAUATWVSH��XH��$�   �E@M�0M�xI���   L��I�͉E�H�M�����wH��PH�UHL�\$0I�ĉ���J��@�E��Ã���!�H��
H�ڄ�HE      DUH��A��L�]��D$ I�KPM�D$L�� L�]�Hcȸ(   )�A�|$  H�M�C��   ���L  H�}H ��   ��   uVH�wHc�H9�|gE��H�G    D��uI�I��L��L���P`H9ظ   E�L��M�u A�uH�e�[^_A\A]A^A_]�@ A�D$N��I��H�wHc�fA�H9�}�H�D6H����U����U�H)�H��L�d$0H�\$(Hc�H�t$ M����� M���_���f�     A�D$L��I��fA��4���f.�     �AH�H��   H�������M�D$A�T$JI�IH)�I�D$L�\$4H�L$(L�L$ L��L�]�I���5� L�]�L)�M��H��H�����������   �����H�}H ������}�@t4����I��A��I�t$LA��A�BH��FfA�AA�D$TfA��v���A�D$T��I��fA��`���������UAWAVAUATWVSH��hH��$�   �EPM�(M�xI���   L��I�̉E�H�M��5��D�sH��PL�@LH��H�UXL�\$0L�E�H��$�   L�]�D��E���J��@�E�@�ƃ���!�@�ƉD$ 襏 �(   L�]�Hc�)ʀ  Hc�M�Suj@����   H�{Hc�H9��  E��H�C    D��uI�E I��L��L���P`H9Ƹ   E�L��M�,$A�\$H�e�[^_A\A]A^A_]�f�     �AH�H��   H����
���L�G�WJI�IH)�H�GL�\$4H�L$(L�L$ L��L�]�I���Y� L�]�L)�M��H��H��@���?���A��   �2���H�}X �'����}�@tlA��H�u���I��A��A�FH��FfA�A�GTfA������ H�D?H����b����U�H)�H��L�t$0H�t$(Hc�H�|$ M���΁ M�����F      ���GT��I��fA�������UWVSH��8H��$�   H��$�   H��$�   H��$�   H��H��A��tpH��H�D$ H)�H��Lc�N�HL�L$(M��I��H���D� D�1�H��H)�H��A)�H��Mc�M��u�*�H��8[^_]�f.�     H��M�H���ra���)���LcH�D$ N�HL�L$(M��I��H���ݏ H)�H���H��8[^_]Ð�����������UAWAVAUATWVSH��   H��$�   )u ���   ���   M�(M�x�E�I���   L�����   H�M`H�M�H�UhL�u�H��H�E����H�{D��L��I��H�ٸ   H��HH��� �CH��0H�t$@%  =  �P  �Z� H�|$ M��H��H�E�H�E�A�-   �t$(H��H�E���� ��,�E���   H�M��
� HcU�H��H�DH����E���L�H)�H��H�D$@H�E�H��H�I���PXLcu�M��M����   �.   M��H��D�u��`��A�T$ H��D�M��  H�M�H)���H�AA�D$Hf���   H�sI9��7  E��H�C    D��uI�E M��H��L���P`L9�   E�H�E`L�(�X(u H�e[^_A\A]A^A_]�D�@Ic�D�E�H��H����d���H)��� D�E�H�t$@�t$(H�M�H�|$ M��H��H�E��Œ �E������A�|$  �N���1�J��   H�������H)��L�t$@��+���h  H�}�A�q��u�   �H��fA�I�FE�L$JL�]�M�D$I�T$H�L$ H�MhH�|$0L��L�\$8H�D$(����u�Lc��u�H�sI9������H�D6H���聲���U�H)�I��H��L�d$@L�t$(Lc�H�t$ M��L����} �u������
� H�}�M��H��G      �t$ A�-   H��H�E�踑 ��,�E������D�@Ic�D�E�H��H�������H)�輧 D�E�M��H��H�t$@�t$ H��H�E��k� �E��p��� �������A��������F<9������V��0��	�����</�����1��t��� L��1�����������UAWAVAUATWVSH��   H��$�   ���   ���   M�(M�x�E�H���   L�uL��H�MpH�MH�Ux�(I���   H��H�E��}��]��H�{D��L��I��H�ٸ   H��HH��[� �CH��@H�t$@%  =  �o  蚦 H�MM��H���m�H�EA�6   H�|$ H�E�H�M�H�D$(�}�H�E��5� ��5�E��   H�M��@� HcUH��H�DH����{���L�H)�H��H�D$@H�E�H��H�I���PXLcuM��M����   �.   M��H��D�u��8\��A�T$ H��D�M��E  H�M�H)���H�AA�D$Hf���   H�sI9��J  E��H�C    D��uI�E M��H��L���P`L9�   E�H�EpL�(�XH�e([^_A\A]A^A_]�fD  D�@Ic�D�E�H��H���蘯��H)��P� D�E�H�t$@M��H�EH�E�H��H�M�H�|$ �m�H�D$(�}���� �E�����     A�|$  �;���1�J��   H����1���H)��L�t$@��+���{  H�}�A�q��u�   �H��fA�I�FE�L$JL�]M�D$I�T$H�L$ H�MxH�|$0L��L�\$8H�D$(����uLc��uH�sI9������H�D6H���褮���U�H)�I��H��L�d$@L�t$(Lc�H�t$ M��L���
z �u�v���f��+� H�}�M��H���m�H�EA�6   H�|$ H�EH��H      H�E��}��̍ ��5�E�����D�@Ic�D�E�H��H�������H)��У D�E�H�t$@M��H�M�H�|$ H���m�H�E�}��y� �E�H�����������A��������F<9������V��0��	�����</�����1��a��� L��1�����������SH��@�Ao H�)D$0L�D$0H��H�L$xH�L$(�L$p�L$ H���PHH��H��@[Ð���SH��@�Ao H�)D$0L�D$0H���L$x�L$(�L$p�L$ H���PH��H��@[Ð����SH��@H��Ao�D$x)L$0L�D$0H���L$p�D$(�L$ H���P8H��H��@[Ð�SH��PH��$�   �Ao �(H��)D$@H�L$0H�H�L$(��$�   L�D$@�|$0�L$ H���P@H��H��P[Ð��SH��@L��  H��AoD�D$xH�@H��)L$0�L$pD�D$(L�D$0L9ЉL$ H��u�+���H��H��@[�f���H��H��@[Ð����SH��@L��  H��AoD�D$xH�@ H��)L$0�L$pD�D$(L�D$0L9ЉL$ H��u�;���H��H��@[�f���H��H��@[Ð����SH��@L�d  H��AoL�D$xH�@(H��)L$0�L$pL�D$(L�D$0L9ЉL$ H��u�����H��H��@[�f���H��H��@[Ð����SH��@L�D  H��AoL�D$xH�@0H��)L$0�L$pL�D$(L�D$0L9ЉL$ H��u�����H��H��@[�f���H��H��@[Ð����VSH��8H��$�   HcL��L��L�D$ L�L$x��L�D$pH�D$(�]v �3H��8[^Ð���UWVSH��XI� I�XA�iH�D$0L�D$0H��L��H��$�   H�\$80ۉ�ᵿ����  H�D$(��$�   A�IH�L$@�D$ �1���H�D$@�n�T$HH�HI      ��H	�H�_H��X[^_]Ð�������������UAWAVAUATWVSH��   H��$�   E�y���   I�8I�XA��I�̋��   A��uRH�M���@��H�}��D$ L�E��t$(H�]������]�H�}��؈�L��I�<$I�\$H�e[^_A\A]A^A_]�fD  I���   L�MxH�M�]���
��@��L�MxD�E�u{Lch@I�qL�X8I9�}{L)�H�D6H����Y���H)�1�L�T$0fE�4BH��H9�u�A��   I�A    A�� tlE��L�]�Hc�uTH�I��L��H���P`L�]�H9�t&A�   �4Lch0I�qL�X(I9�|�E��I�A    uH�M��L��H���P`I9�A��D�É������f�E��L�U�u�H�M��L��H���P`L�U�I9�u�H�Hc�L��H��I���P`H9�A��븐���SH��P��$�   ��$�   �Ao�D$ L�D$@H���D$0�D$(    )L$@����H��H��P[Ð�������SH��`H��$�   �Ao �(H��)D$P�D$(L   H�D$@H�D$0��$�   L�D$P�|$@�D$ �h���H��H��`[Ð��������������SH��@�D$x�Ao �D$(�D$pH��L�D$0)D$0�D$ ����H��H��@[Ð���������SH��@�D$x�Ao �D$(�D$pH��L�D$0)D$0�D$ �����H��H��@[Ð���������SH��@H�D$x�Ao H�D$(�D$pH��L�D$0)D$0�D$ ����H��H��@[Ð�������SH��@H�D$x�Ao H�D$(�D$pH��L�D$0)D$0�D$ ����H��H��@[Ð�������H�99 Ð�������H�AÐ������������/�������������H�Ð�����������SH��01�L�D$/H��1��W H�H��H��0[Ð�������������SH��0H�J      H��H�L$hH�L$(�L$`�L$ H���PH��H��0[Ð���L��   H�H�@L9�u1��f.�     H���������������L�i   H�H�@L9�u1��f.�     H���������������L�I   H�H�@ L9�u�H�����������SH�� H�T$XH���n H��H�� [Ð����1�Ð������������Ð��������������H�Ð�����������SH��01�L�D$/H��1��Z�  H�H��H��0[Ð�������������SH��0H�H��H�L$hH�L$(�L$`�L$ H���PH��H��0[Ð���L��   H�H�@L9�u1��f.�     H���������������L�i   H�H�@L9�u1��f.�     H���������������L�I   H�H�@ L9�u�H�����������SH�� H�T$XH����  H��H�� [Ð����1�Ð������������Ð��������������SH��0H�BH�PL�D$/H���l H��H��0[Ð������������SH��0H�BH�P(L�D$/H���Vl H��H��0[Ð������������SH��0H�BH�P8L�D$/H���&l H��H��0[Ð������������H�Y   H�H�@H9�uH�A�@H�@ H���������������H�9   H�H�@H9�uH�A�@I�@ H���������������H�A�@HÐ������H�A�@IÐ������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P�`k H��H��0[��    H����H��H��0[Ð�SH��0H�H�@(H��H�����H9�u%H�BL�D$/H��H�P(�k H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H�����H9�u%H�BL�D$/H��H�P8��j K      H��H��0[��    H����H��H��0[Ð�SH��0H�BH�PL�D$/H���j H��H��0[Ð������������SH��0H�BH�P(L�D$/H���v�  H��H��0[Ð������������SH��0H�BH�P8L�D$/H���F�  H��H��0[Ð������������H�Y   H�H�@H9�uH�A�@H�@ H���������������H�9   H�H�@H9�uH�A�@J�@ H���������������H�A�@HÐ������H�A�@JÐ������SH��0H�H�@ H��H�����H9�u%H�BL�D$/H��H�P�`i H��H��0[��    H����H��H��0[Ð�SH��0H�H�@(H��H�����H9�u%H�BL�D$/H��H�P(�0�  H��H��0[��    H����H��H��0[Ð�SH��0H�H�@0H��H�����H9�u%H�BL�D$/H��H�P8���  H��H��0[��    H����H��H��0[Ð�H��  H�H�@H9�u1��f.�     H���������������AWAVAUATUWVSH��xH��$�   M�8I�XI�9I��I��M�aH���   H��$�   �`� L��L�|$PH�@H�L$`H�\$XL�L$@H�|$@L�D$PL�d$HH�@H�t$ H�l$(H�D$8H��$�   H�D$0�1  �D$hH�    ����L�|$`H!�H	Ã��@��M����@ �A��uSA�����H��t��u$@8�u�M L��M�>I�^H��x[^_]A\A]A^A_�1�H�WH9Wr�H�H���PH������f�1�I�GI9Gr�I�L���PH����    AD�LD�놐��������AWAVAUATUWVSH��xH��$�   M�8I�XI�9I��I��M�aH���   H��$�   � � L��L�|$PH�@H�L$`H�\$XL�L$@H�|$@L�D$PL�dL      $HH�@ H�t$ H�l$(H�D$8H��$�   H�D$0��  �D$hH�    ����L�|$`H!�H	Ã��@��M����@ �A��uSA�����H��t��u$@8�u�M L��M�>I�^H��x[^_]A\A]A^A_�1�H�WH9Wr�H�H���PH������f�1�I�GI9Gr�I�L���PH����    AD�LD�놐��������AWAVAUATUWVSH��   I�0I�XM�)M�qH��$�   H��H�D$8   L��$  H�D$HH��$  H��$�   �D$0'  L�L$`�D$(    L�D$pH�t$pH�D$@H��$�   H�D$ H�\$xǄ$�       L�l$`L�t$h��  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   D��$�   E�HdE��A������L��$   AH�A�H���@��H����@ �A���|   A�����M��t��u,@8�uA�$H��H�U H�]H�Ĩ   [^_]A\A]A^A_� 1�I�uI9ur�I�E H�T$XL���PHH�T$X�������     A�$�q���fD  1�H�FH9F�t���H�H���PH�    ���AD�HE��V�����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[Ð1�Ð������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[ÐAWAVAUATUWVSH��H�
   I�@I�yI�M�9H�D$0A��H��$�   H��$�   H���   �	� H��$�   I��tH��$�   ��  �   E�A��1�H��=��E1�A�����H�D$(A�����H��@M      ��@ ��(  ��A�����M��t����   1�L;�$�   ��  @����  H��t���  D��A��Hc�A��>9  ��u&I�H�@@H;D$(��   ��*�&  A��>9  �ʍA�<	�  �D� �lAЉ���;�$�   ��   �;�$�   ��   ��A��H�C����H;C�  H��H�CI��A����������     I�GI9G�&���I�D�T$<L���T$8�PH�T$8A����̃��D�T$<�������E1������H�CH9C��   1�������    H�CH;C�  �8��������     D�T$8��A�*   L����D�T$8A����̉�*������    H��$�   ueI��u_��dH��$�   �(H�    ����H#D$0I	�H��$�   H�L�`H��H[^_]A\A]A^A_�H�D�T$8H���PPD�T$8A����������f�H��$�   �� L;�$�   t��q����H�H��D�T$<�T$8�PH�    �T$8A����̃���    D�T$<E�HD�����D  H�D�T$8H���PHA�����D�T$8���t
����������   �����1������������AWAVAUATUWVSH��  L��$�  I�0I�XI�9I��I��M�aI���   H��$�  �� H��$�   Ǆ$�       H�@L�L$`L�D$pH���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$�   H���   H���   H�t$pH�\$xH��$   L��H��$  H��$�   H�|$`H�D$@H�N      �$�   H�D$(H��$�   H�D$ L�l$8H�D$0   L�d$h�  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   H��$�  D��$�   D�A���A��H����D �A��u|A�����H��t��u,A8�u�M L��I�I�^H��  [^_]A\A]A^A_�D  1�H�wH9wr�H�H�T$XH���PHH�T$X������f�     �M �v����    E1�H�FH9F�s���H�H���PH�    ���ED�HE��U����UAWAVAUATWVSH��XH��$�   H�EXH�}P�Ao �Ao	H�M L�mHH���   )E�)M��J� I��H��   H�������H�u�H)�H�E�H��H�E�L�d$ H���'$����t$H�E`�H�E foU�H�e�[^_A\A]A^A_]ËU�H����$��H��A��t�1�E1��%D  I�D�]�L���PD�]�A8�tH��H9�tI�D� �D8�u�C��H��I��H9�u�1�I����   fD  Ic$�   I�L� �?��I��f.�     Ic�I�L� �?��I9�LG�H��I9�w�H�M�H�AH;A�P  H��H�AH���E�����L9�����H�U�H���#���������1��I��C��I9։v4I�<�H�M�HcH��I�D� D�<�E�t	�����   A8�u�H��I9�w�I���/���I�������H�M�H���� Ic$�E�����M�|� A��L���>��H9�H����   �H�U�H���t"�����I����U�H��E�,�\#��A8��0���H�M�H���F� H9��E�����u�H�E@D�0����H�AH;As� �E���H�H�U��PHH�U�����.���H�E�    ��������� H��PP����t���O      ����������������AWAVAUATUWVSH��h  L��$�  I�0I�XI�9I��I��M�aI���   H��$�  轟 H��$�   H�@L�L$`L�D$pH��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$�   H��P  H��$�   H��X  H��$�   H��`  H��$�   H��h  H��$�   H��p  H��$�   H��x  H��$�   H���  H��$�   H���   H��$   H���   H��$  H���   H��$  H���   H��$  H���   Ǆ$�       H��$   H���   H��$(  H���   H��$0  H��   H��$8  H��  H��$@  H��  H��$H  H��  H��   L�l$8H�D$0   H�t$pH��$P  L��H��$X  H��$�   H�D$@H��$�   H�D$(H��$�   H�D$ H�\$xH�|$`L�d$h��  ��$�   H�    ������$�   H!�H��$�   H	Åɉ�H����   H��$�  D��$�   D�A���A��H����D �A��uwA�����H��t��u'A8�u�M L��I�I�^H��h  [^_]A\A]A^A_�1�H�wH9wr�H�H�T$XH���PHH�T$X������f�     �M �{����    E1�H�FH9F�x���H�H���PH�    ���ED�HE��Z����AWAVAUATUWVSH��H  L�=F2��1�H��$�  H��$�  �Ao�AoH���   H��$�  H��H��$�  )�$�   )�$�   �{� H��H�D$X�.� H��I���S:����$�   Ǆ$�       H��$�   H�ƃ��@��H����@ �A���}  ��$�   �H��$�   ��H�P      �t����   1�H9���$�   ��  @����  ����  L�$;E�4$H�oC��59  L����u#I�U L�J@M9���  ����   C��59  ��%��   D�$+C��%9  L����u#I�U L�J@M9���  ����  C��%9  ��Ǆ$�       ��E��   ��O��   ��A��8��  H�=� ��Hc�H���H�AH9A����H��PH�������HǄ$�       �������H��$�   A�<$��$�   H��t	�����   @8��  ��$�   H�$�   �t���f.�     1�H�AH9A�s���H��PH����d���HǄ$�       D���P���H�o�|;A��=9  H��������I�U L�J@M9��  ����   A��=9  ��������     ��uH9�tH��$�  �H��$�  fo�$�    H��H  [^_]A\A]A^A_�@ A��E1�L��A���"���H�AH;A�Q  � @8�������� H������Ǆ$�   ����H��$�   �Y���E1�A��L��A�ф�����f.�     ��$�   ��$�   H��$�   f�     H�}�����    ��$�   H��$�   �����A��=9  ��u#I�M ��L�I@M9���  ���_  A��=9  ��	H��$�   ��  ��$�   ��$�   ��    H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@H�D$8H��$�  L��$�   H��$�  L��$�   H�D$0H��$�   H�D$(H��$�  H�D$ ����H��$�   ��$�   H��$�   ��$�   �����H��$�   H��$�  H�D$8   H�D$Q      HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �&���D��$�   H��$�   ��$�   E��H��$�   ��$�   �'�����$�   H��$�  �G������$�   H��$�   �,��I�U0���B �  H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(
   H��$�  H��$�   H�D$ L��$�   L��$�   �4���H��$�   ��$�   H��$�   ��$�   ��H��$�   ��$�   ��$�   �(�������� H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �i���D��$�   H��$�   ��$�   E��H��$�   ��$�   �j�����$�   H��$�  ���G�P�����$�   H��$�   �l����A��=9  ��u#I�M ��L�I@M9���  ����  A��=9  ��
H��$�   �`����#� H��$�   �����Ǆ$�   ���������fD  H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(   H��$�  H��$�   H�D$ L��$�   L��$�   ����D��$�   H��$�   ��$�   E��H��$�   ��$�   ������$�   H��$�  �G���� H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���  R       H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   )�$�   )�$�   H��$  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ������$�   H��$�   ��$�   ��H��$�   ��$�   �������$�   H��$�  �G�����fD  H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   H��$  H��   H��$  H��  H��$   H��  H��$(  H��  H��$0  H��   )�$�   )�$�   H��$8  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ����D��$�   H��$�   ��$�   E��H��$�   ��$�   �P�����$�   H��$�  �G�9���f�     H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0'  L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �y�����$�   H��$�   ��$�   ��H��$�   ��$�   �|���D��$�   H��$�  E�HdE��A������AH��G�R���f�H��$�   L��L�� I��I�P��%��H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�   ����H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   S      fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(    �)���H�D$XH��$�   fo�$�   fo�$�   H�@H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$   H���   H��$  H���   )�$�   )�$�   H��$  ����f.�     H�D$XH��$�   fo�$�   fo�$�   H�@H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$   H��P  H��$  H��X  H��$  H��`  H��$  H��h  H��$   H��p  H��$(  H��x  H��$0  H���  )�$�   )�$�   H��$8  �;���@ H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@0����@ H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   L��$�   �D$0<   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ����D��$�   H��$�   ��$�   E��H��$�   ��$�   ������$�   H��$�  �����@ H��$�   L��L�� I��I�P���!��H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�   �j���H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@ �)���f���$�   H��$�   H�����I�U0���B�(���H��$�  L��$�   H�D$0   H��$�  L��$�   L�t$@fo�$�   H��$�   L�d$ fo�$�   L��$�   H�L$pH�D$8H��G L��$�   )T      �$�   )�$�   L�L$`H�D$(L�D$h�F���H��$�   H��$�   H��H��$�   ��$�   ��$�   �����$�   ���h�����$�   �$�   �T���H�����A�}8 A���[  A�EfA8�t*��$�   H���f��A�}8 ���P  A�Ed@8�����H��$�  L�t$HH�|$p�D$0   fo�$�   �D$(    L�L$`L�d$ L�D$h)�$�   H��$�  H�D$@H��fo�$�   H�D$8   )�$�   �z���H��$�   L�t$HH��H��$�  L�d$ L�L$`H�D$8   L�D$h�D$0;   H��$�   ��$�   fo�$�   �D$(    )�$�   ��$�   H��$�  fo�$�   )�$�   H�D$@�����H��$�   ��$�   H��$�   ��$�   �����H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   L��$�   �D$0;   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �F���D��$�   H��$�   ��$�   E��H��$�   ��$�   �G�����$�   H��$�  �G�0���H��$�   L��L�� I��I�P�����H��$�   H�|$8fo�$�   fo�$�   )�$�   )�$�   ����@��E1�L��A�������H��$�   ��� H��$�   Ǆ$�   ����fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$0	   �D$(   �����H��$�   ������E1�L��A�щ�������E1�L��A�щ��f���H��PH���tH��$�   ����HǄ$�       1��z����-   L��D$|�3��D�DU      $|�����+   L����������������UAWAVAUATWVSH��XH��$�   H�EX�Ao �Ao	L�}HH�M H���   )E�)M�螈 H��H�EPH��   H����6z��H�]�H)�H�U�H���	��L�t$ ���  �E�1�1�1�H�M�A����� �����H���� �A���  �}��H�M�A��H����D �A����   D8���  D�U�H�M�A���u	H���  H���2  1�E1��I��H��H9�s1H��H92v�I��Lc	O��E81tTH��E��H9�D�	H��H�
r�I9��  H�M�H�AH;A��   H��H�AD�m�H��D���*���f.�     H���f.�     E1�H�AH9A�4���H�D�E��U��PH�U����D�E�����H�E�    E������1�H�AH9A�����H��U��PH�U���������H�E�    D������f.�     H�AH;A��   H��D������D  H�E`�H�E foU�H�e�[^_A\A]A^A_]�H��PPH�M�����H��uH97u�Ic��+UPH��H;MPC�H�U@��H��u�H97t�H9wu��ӋU�H��E1�1��U��H�uPA��H�u ��   @ H�H���PA8�tI��I9�tK���D8�u�E�,�I��H��I9�u�H��H�M�u�E�1�1�����H��PH���tmA���������� H��   �E�����H����gw��M�$�H)�M��H�|$ H��D  IcE I��H��I���"��H�F�M9�u�H�M�������   ����H�E�    A������a����E�H��1�H�M�����������������AWAVAUATUWVSH���   H��$`  H��$x  H��$�  H��$h  H�  V       �Ao H��$@  �Ao)H��H�D$XH��$H  )�$�   )�$�   �Є H9��E     H���/  H��$�   H�D$PH��$�   H�D$HH�,��H�D$`�   f�H�N0���$�   �A �  L�t$HL���{��H����H��P �H��A��H��P D8�t3��$�   L���L��H����H��P�H��A��H��PD8��'  H��$�   H���� Ǆ$�   ����H9��e  �E ���Z  H�T$PH�L$H��������  D�+F��.9  L��E��u*H�L�J@H�n��I9��%  ������B��.9  A��A��%�����L�kL9���  D�[F��9  M��E��u+H�H���H�@@H9��  E����  F��9  E��A��Et
A��O��  L�kL9��,  �[��9  I�߄���  H�H����H�@@H9���  E��tD��9  H�L$Xfo�$�   fo�$�   )�$�   )�$�   趂 �E     �x8 H����  D�`^E��D��$�   ��  D��$�   Ƅ$�    H��$�   H�l$(H��$H  H�D$8H��$p  H��$�   fo�$�   L�L$pfo�$�   L��$�   )�$�   H�D$0H��$`  )\$pH�D$ �o���H��$�   H��$�   H��$�   H��$�   ��$�   ��$�   ������t�M H��$�   I�]H9�H��H��$�   H��$�   H��$�   H��$�   ��$�   ��$�   �����H��$@  fo�$�    H���   [^_]A\A]A^A_�fD  H�CH9��n  D�CH��B�A u�f���A t	H��H9�u�H��$�   A������   ��$�   �H��W      $�   A��H����D �A����   E8��������$�   H��$�   ���u	H����   H�V0���B �����H��$�   H�AH;A��   H��H�AD��$�   D�����A��H����D �A���a���E1�H�AH9A�P���H��PH����A���HǄ$�       E���-����     E1�H�AH9A�:���H��PH����+���HǄ$�       E������H�AH;A��   D� H�V0B�B �C��������fD  H��PPH��$�   �-���D��$�   D��$�   Ƅ$�    �4���H������H�H�@0H;D$`������%   H����A�������@ A��E1�H��A�������E��E1����� A���v����     H��PH����r���HǄ$�       �a���L�\$hA��E1�H����L�\$hA�������f���E1�H����A�������E    �c����E    �W���H�������������������AWAVAUATUWVSH��   H��$   I�8I�XI�)H��I��M�aH���   D��$  D��$   �~ H��$  �    �x8 �  �P^E�툔$�   ��   D��$�   D��$�   Ƅ$�    H��$�   L��H�|$`H�D$8H��$  H�L$pL�L$PH�\$hL�D$`H�l$PL�d$XH�D$0H��$  H�D$(H��$   H�D$ �B����D$xH�    ����L�t$pH!�H	Ã��@��M����@ �A����   A�����H��t����   @8�uH��$  �H��L�6H�^H�Ę   [^_]A\A]A^A_�D��$�   Ƅ$�    ����f�     H��H�D$H���H�D$HH����H�L�B0�%   I9�������%   H��A�X      Љ�����1�I�FI9F�P���I�L���PH����    AD�LD��2���f�1�H�MH9M�4���H�E H���PH��������������������AWAVAUATUWVSH��   H��$   M�0I�XI�9H��I��I�iH���   D��$  D��$   �e| H��$  �    �x8 �  �P^E�䈔$�   ��   D��$�   D��$�   Ƅ$�    H��$�   L��L�t$`H�D$8H��$  H�L$pL�L$PH�\$hL�D$`H�|$PH�l$XH�D$0H��$  H�D$(H��$   H�D$ �"����D$xH�    ����L�t$pH!�H	Ã��A��M����D �A����   �����H��t����   A8�uH��$  �H��L�6H�^H�Ę   [^_]A\A]A^A_�D��$�   Ƅ$�    ����f.�     H��H�D$H�s��H�D$HH����H�L�B0�%   I9�������%   H��A�Љ�����E1�I�FI9F�O���I�L���PH����    ED�LD��1����1�H�OH9O�3���H�H���PH���������������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[ÐH��  H�H�@H9�u1��f.�     H���������������AVAUATUWVSH��   H��$�   �AoI�Y      )M�qI��H��)L$@L��$�   H���   �x foT$@H��H�l$`H�@L�L$`L�t$hH��$�   )T$pL�D$pH�@H�\$ L�l$(H�D$8H��$   H�D$0��  H��$�   H�D$@foD$@fĄ$�   )D$P�D$XH�|$Pfo\$Pf���)\$@��H���� ؉�u_fA�����H���t��u.8�uA�M H�|$@fod$@L��A$$H�Đ   [^_]A\A]A^�H�EH;EsD� f�������     H�GH;Gs6� f����    �    D�HD��z���f�     H�E H���PH�@ H�H���PH�����AVAUATUWVSH��   H��$�   �AoI�)M�qI��H��)L$@L��$�   H���   �w foT$@H��H�l$`H�@L�L$`L�t$hH��$�   )T$pL�D$pH�@ H�\$ L�l$(H�D$8H��$   H�D$0�Y  H��$�   H�D$@foD$@fĄ$�   )D$P�D$XH�|$Pfo\$Pf���)\$@��H���� ؉�u_fA�����H���t��u.8�uA�M H�|$@fod$@L��A$$H�Đ   [^_]A\A]A^�H�EH;EsD� f�������     H�GH;Gs6� f����    �    D�HD��z���f�     H�E H���PH�@ H�H���PH�����AVAUATUWVSH��   �AoI�)M�qL��$  H��$�   I��H�D$8   H�D$HH��$  H��$�   �D$0'  L�L$p�D$(    L��$�   )L$PH�D$@H��$�   H�D$ Ǆ$�       )�$�   H�l$pL�t$x�  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   ��$�   D�Ad�ɍZ      �����H��$   AHЉQf�����H���� ؉�uqfA�����H���t��u.8�uA�M H�|$Pfod$PL��A$$H�İ   [^_]A\A]A^�H�EH;EsV� f�����8�u��fD  A�M �f�     H�GH;Gs6� f����    �    D�HD��h���f�     H�E H���PH�@ H�H���PH�����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[Ð1�Ð������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[ÐAWAVAUATUWVSH��HA�
   I�@I�qI�M�!H�D$0��H��$�   H��$�   H���   �s H��$�   I��tH��$�   A��  �   AD�A��f�����L�d$(@��1�E1�H��A��L��A���   H�|$( D����D ���   H;�$�   D���&  @8��  H��t	E���.  A��H�>A�*   H���W`�PЀ�	�@  C����D�|P�D��A��;�$�   �   D�;�$�   �  �����A��H�CA��A��H;C��   H��H�CH��A�����fA���A��H��@��D ��,���H�CH;C�  � f����    �    HD�E�H�|$( ��D ��	���H�L$(H�AH;A��   � f����    �    E�HEL$(H;�$�   H�L$(�����H��H;�$�   D��uFH��$�   D�8�Yf�H�CH;C��   �f����    HD�����H�H���PP����H��D��H��$�   [      u?H��u9H��$�   E�W�D�H��$�   f�l$0H�t$0H�H�pH��H[^_]A\A]A^A_�H��$�   ���f�H�D�D$>H���PHD�D$>������    H�L$(D�D$?�T$>H��PHD�D$?�T$>�����H�H���PH���,��������������AVAUATUWVSH��   H��$�  �AoI�)M�iI��H��)L$PL��$�  H���   ��o foT$PǄ$�       H��$�   H�@L�L$pL��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$   H�PxH��$  H���   H���   )�$�   H��$  H��H��$  H��$�   H�l$pH�D$@H��$�   H�D$(H��$�   H�D$ H�\$8H�D$0   L�l$x��  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   H��$�  ��$�   �Jf�����H���� ؉�uufA�����H���t��u28�uA�$H�|$Pfod$PL��A&H��   [^_]A\A]A^�D  H�EH;EsV� f������f.�     A�$�f�     H�GH;Gs6� f����    �    D�HD��d���f�     H�E H���PH�@ H�H���PH�����UAWAVAUATWVSH��hH��$�   H�EhL�e`�Ao �Ao	H�M0H�]XH���   )E�)M���m I��J��   H����&_��H�U�H)�H�E�H�U�H�E�L�|$ H��������t$H�Ep�H�E0foU�H�e�[^_\      A\A]A^A_]��U�H�M��A���M���t�1�E1�� I�L���P0f9�tH��I9�tH���f9�u�C�4�H��I��I9�u�1�I����   Ic7A�   H���	��I��Kc�H���	��I9�LG�I��M9�r�H�M�H�AH;A�l  H��H�AH�������L9�f�U�����H�U�H�M������������L�?1���I��C��I9�A��v2Ic4�H�M�H��H��B�4�E�t
f�����   f9�u�H��I9�w�I���3���I�������H�M�H����� �����f�E�IcH�4�A��H�����H9�I��sQA����� L�}�H�U�L���������V����U�L���~����f9��=���H�M�H���� L9�fD�u�r�I9�����H�EPD�(���� H�AH;As� f����.���H�E�    �!���H�L�M�H�U��PHL�M�H�U���@ H��PP���������AVAUATUWVSH��p  H��$�  �AoI�)M�iI��H��)L$PL��$�  H���   �lj H��$�   H�@L�L$pL��$�   H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$�   H��P  H��$�   H��X  H��$�   H��`  H��$�   H��h  H��$�   H��p  H��$�   H��x  H��$   H���  H��$  H���   H��$  H���   H��$  H���   H��$   H���   H��$(  H���   foT$PǄ$�       H��$0  H���   H��$8  H���   H��$@  H��   H��$H  H��  H��$P  H��  H��$X  H��  H��   H�\$8H�D$0]         )�$�   H��$`  H��H��$h  H��$�   H�D$@H��$�   H�D$(H��$�   H�D$ H�l$pL�l$x�  H��$�   ��$�   H�D$PfoD$PfĄ$�   )D$`fo\$`��H�|$`)\$P�D$h��   H��$�  ��$�   �Jf�����H���� ؉�upfA�����H���t��u-8�uA�$H�|$Pfod$PL��A&H��p  [^_]A\A]A^�H�EH;EsV� f������f.�     A�$�f�     H�GH;Gs6� f����    �    D�HD��i���f�     H�E H���PH�@ H�H���PH�����AWAVAUATUWVSH��H  L�5�� E1�H��$�  H��$�  �Ao�AoH���   H��$�  H��H��$�  )�$�   )�$�   ��f H��H�D$X�g H��H�������$�   Ǆ$�       H��$�   I��H��$�   H�D$`f���@��H����@ ����n  f��$�   �H��$�   ��H���� Љ���   @8׋�$�   ��   M9���   ����   H�K�,$E1�H��L�,.A�U I�|$�P`<%uGH�E1�H���T.�P`Ǆ$�       <E�  <O�  ��A<8�I  ��Ic�L���@ H��$�   A�m ��$�   H��t
f����=  f9��c  ��$�   I����$�   �����H�AH;A�   � 1�f��������ꋄ$�   HǄ$�       @8�������uM9�tH��$�  �H��$�  fo�$�    H��H  [^_]A\A]A^A_�@ H�AH;A��  � 1�f����u���HǄ$�       ���b���H�I�|$E1�H���T.�P`��^      ���D  ��$�   H�L$`�N���E1�H����H��P`<	�"  ��$�   ��$�   �    L�gH��$�   �����H�AH;A��  � f�����  f9�H��$�   ����� �� �����I��H��$�   f��$�   ���������f�     H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@H�D$8@ H��$�  L��$�   H��$�  L��$�   H�D$0H��$�   H�D$(H��$�  H�D$ �L���H��$�   ��$�   H��$�   f��$�   ������    H�D$XH��$�   fo�$�   fo�$�   H�@H�PXH��$�   H�P`H��$�   H�PhH��$�   H�PpH��$�   H�PxH��$   H���   H��$  H���   )�$�   )�$�   H��$  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ �)���H��$�   ��$�   H��$�   ��$�   f��$�   ���������$�   H��$�  �A���� H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$   H���   H��$  H���   H��$  H��   H��$  H��  H��$   H��  H��$(  H��  H��$0  H��   )�$�   )�$�   H��$8  H��$�   H��$�  H�D$0   H�D$@H��$�  L��$�   L��$�   H�D$8H��$�   H�D$(H��$�   H�D$ ����H��$�   ��$�   H��$�   ��$�   _      f��$�   ���@�����$�   H��$�  �A�)���f�     H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0'  L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �)�����$�   H��$�   ��$�   ��H��$�   f��$�   �j�����$�   D�Ad�ɍ�����H��$�  AH��A�C��� H�L�U� H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   H�l$8����H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(    H��$�  H��$�   H�D$ L��$�   L��$�   �������$�   H��$�   ��$�   ��H��$�   f��$�   �7�����$�   H��$�  �A� ���H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(   �.���H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0;   L��$�   fo�$�   �D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �����D��$�   H��$�   ��$�   E��H��$�   f��$�   ������$�   H��$�  �A�����H�L�
� H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   �����H��$�   H��$�  H�D$8   H�D$HH��$�  L��$�   H��$�   �D$0<   fo�$�   �`      D$(    L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   ����D��$�   H��$�   ��$�   E��H��$�   f��$�   �������$�   H��$�  ������f�H�L��� H��H��$�   I�P�I���PXH��$�   fo�$�   fo�$�   )�$�   )�$�   ����f�H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@ H�D$8�������$�   H�L$`�M���L��   H��D��A�Q�������H��$�  L��$�   H�D$0   H��$�  H��$�   M��fo�$�   L��$�   H�l$@fo�$�   H��$�   L�l$ H�D$8H�n L��$�   H�L$p)�$�   )�$�   H�D$(L�D$h����H��$�   H��$�   H�L$`H��$�   ��$�   f��$�   ������$�   ���@�����$�   �$�   �,���H�L$`�B����-   H��f�D$~H��PPf9D$~t0��$�   H�L$`�����+   H��f�D$~H��PPf9D$~�����H��$�  M��H�l$Hfo�$�   �D$0   L�D$hL�l$ H��$�  )�$�   H�L$pH�D$@fo�$�   �D$(    H�D$8   )�$�   �����H��$�   H�l$HM��H��$�  L�l$ L�D$hH�D$8   H�L$p�D$0;   H��$�   ��$�   fo�$�   �D$(    )�$�   f��$�   H��$�  fo�$�   )�$�   H�D$@�p���H��$�   ��$�   H��$�   f��$�   ����H�D$XH��$�   fo�$�   fo�$�   H�@H���   H��$�   H���   H��$�   H���   H��$�   H���   H��$a      �   H���   H��$   H���   H��$  H���   )�$�   )�$�   H��$  �����f.�     H�D$XH��$�   fo�$�   fo�$�   H�@H��(  H��$�   H��0  H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$   H��P  H��$  H��X  H��$  H��`  H��$  H��h  H��$   H��p  H��$(  H��x  H��$0  H���  )�$�   )�$�   H��$8  �[���@ H�D$XH��$�   fo�$�   fo�$�   )�$�   H�@)�$�   H�@0H�D$8����H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�   H�D$@H��$�   H�D$ )�$�   �����H��$�   ��$�   H��$�   ��$�   f��$�   ���)�����$�   H��$�  �A����f���$�   H�L$`����L��    H��D��A�Q���  H��$�   �D$0   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$(
   H��$�  H��$�   H�D$ L��$�   L��$�   �����H��$�   D��$�   H��$�   ��$�   E��f��$�   ��$�   �#����������$�   H�L$`�,���E1�H����H��P`<
�����H��$�   �� A����������fD��$�   �����H��$�   H��$�  H�D$8   H�D$HH��$�  H��$�   �D$0   L��$�   fo�$�   �D$(   L��$�   fo�$�   )�$�  b       H�D$@H��$�   H�D$ )�$�   �����D��$�   H��$�   ��$�   E��H��$�   f��$�   ������$�   H��$�  ���A�����H��PH�����f�H��PH�f���D  HǄ$�       1�����H��$�   A�����躴 H��$�   fD��$�   fo�$�   H�D$HH��$�  H��$�   fo�$�   )�$�   H�D$8   )�$�   H�D$@�D$0	   �D$(   �����H��PH�f�������UAWAVAUATWVSH��XH��$�   H�EX�Ao �Ao	L�uHH�M H���   )E�)M��^T I��H�EPH��   H����E��H�]�H)�H�U�H���3���L�l$ ���  H�M�1�1�1��E�A�����f�f���A��H����D ����G  f�}��H�M���H���� �A����   A8���   �E�H�M�f���u	H���:  H����   L�61�E1��fD  I��H��H9�s4H��H91v�M�D� McO��fC9tHH��E�T� H9�E�L��L�r�I9�tkH�M�H�AH;A��   H��H�AfD�}�H��D������H���f�     H�AH;A��  � 1�f����)���D��H�E�    A8�����H����   H97��   H�E`�H�E foU�H�e�[^_A\A]A^A_]��     H�AH;A��  � E1�f��������H�E�    A������f�H�AH;A�c  � f��������H�E�    �����     H��PPH�M�����H���[���H97t
H9w�L���IcM ��+UPH��H;MPC�H�U@��5����U�H��E1�1�����H�uP��H�u%��   f�     I�L���P0f9�tI�c      �I9�tK���f9�u�E�d� I��H��I9�u�1�1�H��H�M��~����5� �����f�E�H��   H�����B��M�d� H)�M��H�|$ H���     IcI��H��I�������H�F�M9�u�H�M��   ����H�D�E��PHD�E�����H��U��PH�U��p���H��PH����H�M�H��1������������AWAVAUATUWVSH���   H��$P  H��$h  H��$p  L��$X  H�   �Ao H��$0  �Ao)H��H�D$PH��$8  )�$�   )�$�   �P H9�A�$    H���z  H��$�   L��$�   H�D$HL��$�   �   f.�     H��    H��D��P���|  ��$�   L�������H����H��P@�H�ى�H��P@f9�t3��$�   L������H����H��P0�H�ى�H��P0f9���  H��$�   H���S� �����f��$�   H9���  E�$E����  L��L���������8  H�E1�H����P`<%�&���H�~H9��!  H�E1�H���V�P`<EA���  <O�	  H�L$Pfo�$�   fo�$�   )�$�   )�$�   �
O A�$    �%   L� H��A�PPf��$�   fE��1�fD��$�   f��$�   H�L$HL�L$`L�d$(H��$�   H��$8  H�D$8H��$`  L�D$pfo�$�   fo�$�   )D$pH�D$0H��$P  )L$`H�D$ �O���H��$�   H��$�   H��$�   H��$�   ��$�   f��$�   �:�����tA�$H��$�   H�wH9�H��H�D$pH��$�   H��$�   H�D$x�D$xf��$�   �U���H��$0  fo�$�    H���  d       [^_]A\A]A^A_�f.�     H��    H��D��P��t	H��H9�u���$�   �����H��$�   �   �    f��$�   �H��$�   ��H���� �A����   A8������H��$�   D��$�   H��tfA�����   H��    H���P���u���H��$�   H�AH;A��   H��H�Af��$�   ��f���A��H����D ����Z���H�AH;A�\  � E1�f����<���HǄ$�       A���(����     H�AH;A�  � 1�f����(���HǄ$�       D������H�AH;A�  D� fA����!���HǄ$�       �����H��PPH��$�   �0���H�~H9���   H�E1�H���V�P`H�L$Pfo�$�   f��fo�$�   )�$�   )�$�   ��K A�$    �%   L� H��A�PPE��f��$�   tofE��1�f��$�   fD��$�   f��$�   ������    H�D�D$_�PHD�D$_�����f.�     H��T$_�PH�T$_����H��PHD�������A���Z���A�$   �F���A�$   �9��������������AWAVAUATUWVSH��   )�$�   H��$   �Ao8I�)M�iI��I��H��$(  )|$@H���   ��$8  D��$@  ��J �%   L� �    H��f��A�PPE��f��$�   �  1�f��$�   f��$�   H��$�   H�t$ L��H�D$8H��$0  L�L$`H��$�   H�|$(L�D$p)|$pH�l$`H�D$0L�l$h����H��$�   H�D$@foD$@fĄ$�   )D$P�D$XL�t$PfoL$Pf���)L$@��M���� ؉���   fA�����H��e      �t��u98�u�L�t$@(�$�   L��foT$@A$H�ĸ   [^_]A\A]A^A_� H�EH;Esf� f������f.�     fE��1�f��$�   fD��$�   f��$�   �����I�FI;Fs1� f����    �    D�LD��H���@ H�E H���PH�@ I�L���PH�ǐ����AWAVAUATUWVSH��   H��$  �AoI�)M�iI��I��)L$@H��$  H���   ��$(  D��$0  �H �%   L� �    H��f��A�PPE��f��$�   �  1�f��$�   f��$�   H��$�   foT$@H�t$ L��H�D$8H��$   L�L$`H��$�   H�|$(L�D$p)T$pH�l$`H�D$0L�l$h����H��$�   H�D$@foD$@fĄ$�   )D$P�D$XL�t$Pfo\$Pf���)\$@��M���� ؉���   fA�����H���t��u.8�u�L�t$@fod$@L��A$$H�Ĩ   [^_]A\A]A^A_�H�EH;Esc� f�������    fE��1�f��$�   fD��$�   f��$�   �����I�FI;Fs1� f����    �    D�LD��V���@ H�E H���PH�@ I�L���PH�ǐ����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[ÐSH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[ÐAWAVAUATf      UWVSH��   ��$�   M�xH��$   L��$  L��$�   I��M�(�D$OH��$�   H��$�   D�|$@H���   �.E L9�D�L$@H����  H�D$pL��$�   M��M��H�D$PH�D$`E��H�D$XH�����H�D$@�2f�     E��uI�F(I;F0���  �I�F(I9�H���A  �+H�{��.9  H���uH�H�@@H;D$@�_  ��t���.9  ��<%u�I9���   �k��.9  H���u$H�H�@@H;D$@�P  ���  ��.9  �р�Et	��O��   H�{I9���   �k����.9  H�����u!H�@��H�@@H;D$@�  ��t��.9  H��$�   E��H��H��$�   L��$�   L�D$XH� H�@�T$0�T$OL�t$`L�l$h�\$8H��H�L$(H�L$P�T$ H��$�   ��D�l$xI9�L�t$pE�������E��M��M��H��$�   E��L�(L�xH�Ĉ   [^_]A\A]A^A_��    1�1��N����    @��E1�H���Љ�����I�L���Ph���A���E����     H��@��E1��Љ�����H��E1����Љ�����������������SH��P�Ao H�)D$@L�D$@H����$�   �L$8��$�   �L$0H��$�   H�L$(��$�   �L$ H���PH��H��P[Ð�����AWAVAUATUWVSH���   M� M�hD��$@  ��$H  I���   H��H���5B H��H���jA �{8 I����   �C^@��D$<��   @�l$=D�t$>�D$? H��$8  H�t$@A��   L��L�L$<H��H��H�D$ �����H����������!�%����t��D�������  D�H�S��HD� �H��H)�E��uI�g      $I��H��L���P`H9ø   E�H��L�'@�oH���   [^_]A\A]A^A_�f.�     D�t$=�D$> �D����H������H�H�����L�@0�%   I9������%   H��A�������������������AWAVAUATUWVSH��   H��$   L��$  M�xI�8H��$�   I���   I��D��$�   L��$�   �A L9�D��H���
  H�D$pH�D$HH�D$`H�D$PA��M���D$X�5@��u$H�O(H;O0��(  f�H��H�O(f���@��M9�L����   H�L�{E1�H����P`<%u�M9���   H�E1�H���S�P`D��A��E��   1�A��O��   I�E A��I��L�D$PL��H�L$HH�@H�|$`H��$�   L�t$h�T$8L��D�L$0L��$�   H�|$(�|$X�|$ ��D�t$xM9�H�|$pD���O���M��H��$�   A��H�8L�xH�Ĉ   [^_]A\A]A^A_�L�{D�L$_M9�t�H�E1�H���S�P`�T$_D���D��� ��H�H���Ph��������������������SH��P�Ao H�)D$@L�D$@H����$�   �L$8��$�   �L$0H��$�   H�L$(��$�   �L$ H���PH��H��P[Ð�����AVAUATUWVSH��@  I�(M�`��$�  ��$�  M���   H��L����> L��f��I���> �%   L��I��I��PP@��f�D$8u1�f�\$:f�T$<H��$�  H�|$@L��A��   L�L$8H��E��H�D$ �g���H�������E��Hc�uH�E I��H��H���P`H9ø   DE�H��H�.D�nH��@  [^_]A\A]A^�f@��1�f�\$<f�|$:f�D$>�r�������H��� Ð��������AÐ������������A ��Ðh      ���������A ���Ð������H���   Ð��������A ��Ð�������VSH��(���    H��t���   H��([^�H���   H��tQ�~8 t�FY���   ƃ�   H��([^�fD  H���X���H�H�����L�@0�    I9�tƺ    H��A���� ���������������A ����Ð������H���   Ð�������VSH��(H���   H�ۉ�tI�{8 t���D39H��([^��    H�������H�H�����L�@0��I9�t�@��H��H��([^I��� ��������������WVSH�� H���   H��D��A��tM����;9  ��u%H�H�����H�@@H9�uD8Ɖ�tD��;9  D��H�� [^_�D����H����A����� ������A Ð������������    �A HD�Ð��A ��Ð��������A ��Ð��������AÐ������������A ��Ð���������A ���Ð������H���   Ð��������A ��Ð�������SH�� ���    H��t���   H�� [�f�H���   H��tH��    �PPƃ�   f���   H�� [��� �����������������A ����Ð������H���   Ð�������H��(H���   H��tH���H�@PH��(H���j ����������H��(H���   H��tH���E��H�@`H��(H���6 �������A Ð������������    �A HD�Ð��A ��Ð��������A ��Ð�������H��� Ð�������AWAVAUATUWVSH��   H��$   �Ao �Ao	H���   H��$   H��)�$�   )L$p��9 H��$�   H��H�D$P袍���D$n H��H�~@ H�@dHi      �D$@t
H�~P �D$nH��$�   1�1�I��H�D$8���  �~  H��$�   tH��$�   �    ��  L��$�   1�1���  H�L$8�    H��$�   �_�  H�FeE1�E1��D$o H�D$0�F`1��D$h    H�D$H    ��$�   H��$�   H�D$XH�D$XB�<0��  B�0H�=m� Hc�H���A�   I����  H�|$H��D!���8  �|$o �=  L�n8L�d$p�   A�����H��$�   �H��H�AD��$�   H��L��H���p���H;|$H�  <�  ��$�   H���N���A8D= �E  H��$�   H�AH;Ar�H��PP�f�     ��$�   L��$�   H��$�   �U�    H�=�� H+D$@H�L$8H���S�  ��H��$�   H�AH;A�z  H��H�AǄ$�   ������������@��H��@��@ ���  �|$x�H�L$p��H��@��@ ���  @8���  ��$�   H��$�   ���u	H����  H�L$0@��A�
   �����H���;���@8~!A��E���  �F ���   @8~"��  E���P  ���P  ��L���h�  1������H��$   �@uRH�|$H@��E����@�u=A���d  A��A�   �{  ��$�   <t<�}  �|$n �r  @ H�F0L�d$pE1�H��$�   H�D$`�>D  ��$�   H���a���H�V(B8*��  H��$�   �F� Ǆ$�   ����I��L��H���,�����L;l$`����@ �u�L;l$`�O  A�   ��   @ L�d$pH��$�   L��H����������  E1�I������L�d$p�����H��$�   �7H�T$P�j      �H�R0�B toH��$�   H�AH;A�7  H��H�A��$�   L��H���}�����u;��$�   H��$�   ���u�H��t�H�AH;A�"  H�T$PD� H�R0B�B u�D���A�F���_���@���V���H�D$XI��B�<0����1�������    H�~@ ��  H�~P L�d$pH��$�   �M  �|$nA��A���1�H�AH9A�$���H��PH�������HǄ$�       ������1�H�AH9A����H��PH1҃�������H�D$p    �������H�AH;A��  �8�����fD  H��PPH��$�   �{����FX����  �\$hA�   1��A���A��H��$�   H�x� �����L�d$pH��$�   H��$(  �L��H��������tH��$(  �H��$   fo�$�   H��$�   H��H��$�   H�H��	�  H��$�   H��H�H����  H��$   H�ĸ   [^_]A\A]A^A_�f�     L�nH�����    L�d$pH��$�   L��H���H��������'  H�~P ��   H�~@ �K���1�A�   �D$o�����fD  ��$�   H������H�|$P��H�W0�B ����H��$�   �ވ Ǆ$�   ����A�   ������     M�������H��$   �@�D$`%   A��@���^���fD  L��H��腳��������  H�~@ �����H�~P ������8���H��PP�����D  H;|$H�G���H��$�   H�x���   �|$o �  H��$�   H�x� t=�D$h��E��H��$�   H��E��j�  H�VI��H�N� ��uH��$(  �E��uvH�T$8H��$0  �$�  L�d$k      pH��$�   ����f�H��PH������G���HǄ$�       ������1���E1�fD  H��$�   A�   H�x� �)����W���f�9^X�L����|���f�H�L$8E1��0   �.g��H������H�����  H�L$8I��1��|�  �������$�   H������H�V88�����H�F@H��$�   H�D$H�� Ǆ$�   ����A�   ������$�   H�������H�VH8�:���H�FPH��$�   H�D$H蟆 A�   �D$oǄ$�   �����L���@ E���l���H��$�   H�x��2��������|$n@���������$�   �������$�   �&�������H��PH����b���HǄ$�       �Q���H�|$8H�����  H��$�   �80�����H����  �D$ -   E1�1�H��A�   ��  H��$�   �@���������E������E1�����H��$�   H�@�H���k���H��$�   H��H��$�   H��H�H����  H��$�   H��H�H����  H����$��H��$�   H���א�������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H���   H��$   H��)�$�   )L$p��. H��$�   H��H�D$P�����D$n H��H�~@ H�@dH�D$@t
H�~P �D$nH��$�   1�1�I��H�D$8���  �~  H��$�   tH��$�   �    ��  L��$�   1�1���  H�L$8�    H��$�   ��  H�FeE1�E1��D$o H�D$0�F`1��D$h    H�D$H    ��$�   H��$�   H�D$XH�D$XB�<0��  B�0H�=y� Hc�H���A�   I����  H�|$H��D!���H  �|$o �M  L�n8Ll      �d$p�   A�����H��$�   �H��H�AD��$�   H��L��H��萮��H;|$H��  <��  ��$�   H���n���A8D= �U  H��$�   H�AH;Ar�H��PP�f�     ��$�   H��$�   H��$�   �U�    H�=�� H+D$@H�L$8H���s�  ��H��$�   H�AH;A��  H��H�AǄ$�   ������������@��H��A��A ���  �|$x�H�L$p��H��A��A ���  @8���  ��$�   H��$�   ���u	H����  H�L$0@��A�
   ����H���;���@8~!A��E���  �F ���  @8~"�  E���`  ���`  ��H����  1������H��$   �@uRH�|$H@��E����@�u=A���t  A��A�   �{  ��$�   <t<�}  �|$n �r  @ H�F0L�d$pE1�H��$�   H�D$`�D  H��H�AǄ$�   ����I��L��H���n�����L;l$`����@ ���  ��$�   H���I���H�V(B8*��  H��$�   H�AH;Ar�H��PP뙐L�d$pH��$�   L��H����������  E1�I������L�d$p�����H��$�   �7H�T$P��H�R0�B toH��$�   H�AH;A�  H��H�A��$�   L��H��蝫����u;��$�   H��$�   ���u�H��t�H�AH;A�2  H�T$PD� H�R0B�B u�D���A�F���_���@���V���H�D$XI��B�<0����1�A�   ��@ H�~@ ��  H�~P L�d$pH��$�   �-  �|$nA��A���1�H�AH9A�$���H��PH�������m      HǄ$�       D������1�H�AH9A����H��PH1҃�������H�D$p    D�������f.�     H�AH;A��  �8�����f.�     H��PPH��$�   �k����FX���{  �\$hA�   1��1���A��H��$�   H�x� �����L�d$pH��$�   H��$(  �L��H���������tH��$(  �H��$   fo�$�   H��$�   H��H��$�   H�H���  H��$�   H��H�H���  H��$   H�ĸ   [^_]A\A]A^A_�f�     L�nH�����    L�d$pH��$�   L��H���X��������*  H�~P uwH�~@ �?���1�A�   �D$o�����f.�     ��$�   H������H�|$P��H�W0�B �����H��$�   ��} Ǆ$�   ����A�   ������     L��H���Ũ��������  H�~@ �����H�~P ������d���H��PP�����D  H;|$H�w���H��$�   H�x��  �|$o �G  H��$�   H�x� t=�D$h��E��H��$�   H��E���  H�VI��H�N�� ��uH��$(  �E����   H�T$8H��$0  �`�  L�d$pH��$�   �����H��PH������e���HǄ$�       ������O���E1�@ H��$�   A�   H�x� �I�������f�L;l$`�i���M���~���H��$   �@�D$`%   A��@������9^X�G����K���H�L$8E1��0   �;\��H�������H����}  H�L$8I��1���  ������$�   H������H�V88�����H�F@H��$�   H�D$H��{ Ǆ$�   ����A�   ������$� n        H���Χ��H�VH8����H�FPH��$�   H�D$H�{ A�   �D$oǄ$�   �����9����E���l���H��$�   H�x����������|$n@���������$�   �������$�   ��������H��PH����R���HǄ$�       �A���H�|$8H�����  H��$�   �80�����H�����  �D$ -   E1�1�H��A�   ��  H��$�   �@������d���E������E1�����H��$�   H�@�H���n���H��$�   H��H��$�   H��H�H����  H��$�   H��H�H����  H������H��$�   H���א�������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����AWAVAUATUWVSH��   )�$�   H��$  �Ao9I�0I�XH��I��D��$   H���   �# L�l$w1�1�M��I���S�  E��H�t$PL��H�D$xH�D$xH�D$0H��$  H�L$`H�\$XL�L$@)|$@L�D$PH�l$ H�D$(��   ����H�D$`H�T$hH�L$xH�D$`H��H�T$h�D$hH�    ����H�i�H!�H	�H��tjH��$  E1�H����  H��$  L�8A�G�����   A�F8L�d$x<t����   I�H�����H�@8H9���   L��I��L��赿��H�L$xH�7�����H�_��A���~+(�$�   H��H�Ę   [^_]A\A]A^A_����������f�o      H��L���$�  ��f�H��$  ���  H��$  L�8�S��� L�������Y��� M��L��L��M�,��H�L$x�g���H��H�D$xL��H�H����  H�����������������AVAUATUWVSH��   )�$�   I�M�h�Ao9D��$�   H�l$xH��H��L��$   1�1�I���T�  H�L$`H�\$PH��H�D$pH�D$pE��H�D$0H��$�   L�L$@L�l$XL�D$P)|$@L�d$(H�D$ ��   ����H�    ����H�D$`H�T$hL!�H��H�D$`H�T$h�D$hH	��� H�L$pI��M��H�D$xH��$  �7� H�L$pH������H�w��A���~-(�$�   H��H�Đ   [^_]A\A]A^������r���fD  H��H���t�  ��H��H�D$pH��H�H��n�  H�����������AWAVAUATUWVSH��   H��$   �Ao �Ao	H���   H��$   H��)�$�   )L$p�  H��$�   H��H�D$P��u���D$j H��H�{@ H�@dH�D$@t
H�{P �D$jH��$�   1�1�I��H�D$8��  �{  H��$�   tH��$�   �    �g�  L��$�   1�1��v�  H�L$8�    H��$�   �?�  H�CfE1�E1��D$k H�D$0�C`1��D$l    H�D$H    ��$�   H��$�   H�D$XH�D$XB�<0��  B�0H�=ݠ Hc�H���A�   I���7  H�|$H��D!����  �|$k ��  L�k8L�d$p�   A�����H��$�   �7fA9D} �*  H��$�   H�AH;A�<  H��H�AfD��$�   H��L��H���}���<�  H;|$H�  H��$�   ��$�   H��t�f���u�H�AH;A�@  � f����p      u���HǄ$�       �d�����$�   L��$�   H��$�   f���@��H��@��@ ���  f�|$x�H�L$p��H��@��@ ���  @8��  H��$�   ��$�   H��t
f�����  H�T$0H�Kz@ f9��  H��H9�u�f9C"��D���  D�k E����  f9C$��  E����  ����  @��L���i�  1�H��$�   H�AH;A��  H��H�A����������f��$�   ����H��$   �@uNH�|$H@��E����@�u9A����  A��A�   �j  ��$�   <t<�l  �|$j �a  H�C0L�d$pE1�H��$�   H�D$`�H��H�AA�����I��fD��$�   L��H���u�����L;l$`����@ ���  ��$�   H������H�S(fB9j��  H��$�   H�AH;Ar�H��PP�H�{@ ��  H�{P L�d$pH��$�   �g  �|$jA��A���  L�d$pH��$�   L��H���ڝ������  E1�I�������L�d$p�����H��$�   �?�H�L$P�    H��P���'  H��$�   H�AH;A�  H��H�Af��$�   L��H���g�������  H��$�   D��$�   H��t�fA���u�H�AH;A��  D� fA����u���HǄ$�       �d���@ H�I� H+T$@H�L$8H� H�����  �������     H�AH;A�  � 1�f��������H�D$p    ��@8������A�   H��$�   H�x� �%  L�d$pH��$�   H��$(  �L��H���s�����tH��$(  �H��$   fo�$�   H��$�   H��H��$�q         H�H��D�  H��$�   H��H�H��0�  H��$   H�ĸ   [^_]A\A]A^A_�@ H�AH;A�F  � 1�f��������HǄ$�       �������H�AH;A�!  � f�������HǄ$�       �����@ H��PPH��$�   �d����KX���  �t$lA�   1��*���D���A�F���b���@���Y���H�D$XI��B�<0� ���1�A�   ��L�kH�U���L�d$pH��$�   L��H�����������  H�{P uiH�{@ �����1�A�   �D$k���$�   H��蛛��H�L$PD���    L�	A�Q��A�������H��$�   �Nx �����f��$�   ����L��H��葚��������  H�{@ �y���H�{P �n����r���H��PP�����H��PP�����H;|$H�����H��$�   H�x���   �|$k �7  H��$�   H�x� t>�D$l@��E��H��$�   H��E���  H�SI��H�K�O� ��uH��$(  �E��uzH�T$8H��$0  �ٿ  L�d$pH��$�   �9���H��PH�����H��PH����H��PH�����L;l$`�L���M�������H��$   �@�D$`%   A��@�������9sX������x���H�|$8E1��0   H����L��H�������H��$�   H���A�    H��L�B�I�P�HD�L9�LF�1����  �������$�   H��豙��H�S8f9�����H�C@H��$�   H�D$H�nv A�����A�   fD��$�   �I�����$�   H���d���H�SHf9����H�CPH��$�   H�D$H�!v A�����A�   �D$kfD��$�   �����f�E�������H��$�   H�x��r      ��������H��PHD��� ����|$j@���l�����$�   �^�����$�   ������K���H��PH����H��$�   �P���ye�80������@���yIH�L$8A�   E1�1��D$ -   �J�  H��$�   �@������y���E1������A�������E�������H�L$8�D�  �H�L$8�8�  H��$�   �E1�����H��$�   H��H��$�   H��H�H��W�  H��$�   H��H�H��C�  H���k
��H��$�   H���א�������������AWAVAUATUWVSH��   H��$   �Ao �Ao	H���   H��$   H��)�$�   )L$p�� H��$�   H��H�D$P�k���D$j H��H�{@ H�@dH�D$@t
H�{P �D$jH��$�   1�1�I��H�D$8�g�  �{  H��$�   tH��$�   �    �'�  L��$�   1�1��6�  H�L$8�    H��$�   ���  H�CfE1�E1��D$k H�D$0�C`1��D$l    H�D$H    ��$�   H��$�   H�D$XH�D$XB�<0��  B�0H�=�� Hc�H���A�   I���7  H�|$H��D!����  �|$k ��  L�k8L�d$p�   A�����H��$�   �7fA9D} �*  H��$�   H�AH;A�<  H��H�AfD��$�   H��L��H���=���<�  H;|$H�  H��$�   ��$�   H��t�f���u�H�AH;A�@  � f����u���HǄ$�       �d�����$�   L��$�   H��$�   f���@��H��@��@ ���  f�|$x�H�L$p��H��@��@ ���  @8��  H��$�   ��$�   H��t
f�����  H�T$0H�Kz@ f9��  H��H9�s      u�f9C"��D���  D�k E����  f9C$��  E����  ����  @��L���)�  1�H��$�   H�AH;A��  H��H�A����������f��$�   ����H��$   �@uNH�|$H@��E����@�u9A����  A��A�   �j  ��$�   <t<�l  �|$j �a  H�C0L�d$pE1�H��$�   H�D$`�H��H�AA�����I��fD��$�   L��H���5�����L;l$`����@ ���  ��$�   H���ϓ��H�S(fB9j��  H��$�   H�AH;Ar�H��PP�H�{@ ��  H�{P L�d$pH��$�   �g  �|$jA��A���  L�d$pH��$�   L��H��蚒������  E1�I�������L�d$p�����H��$�   �?�H�L$P�    H��P���'  H��$�   H�AH;A�  H��H�Af��$�   L��H���'�������  H��$�   D��$�   H��t�fA���u�H�AH;A��  D� fA����u���HǄ$�       �d���@ H�	� H+T$@H�L$8H� H������  �������     H�AH;A�  � 1�f��������H�D$p    ��@8������A�   H��$�   H�x� �%  L�d$pH��$�   H��$(  �L��H���3�����tH��$(  �H��$   fo�$�   H��$�   H��H��$�   H�H���  H��$�   H��H�H���  H��$   H�ĸ   [^_]A\A]A^A_�@ H�AH;A�F  � 1�f��������HǄ$�       �������H�AH;A�!  � f�������HǄ$�       �����@ H��PPH�t      �$�   �d����KX���  �t$lA�   1��*���D���A�F���b���@���Y���H�D$XI��B�<0� ���1�A�   ��L�kH�U���L�d$pH��$�   L��H���֏�������  H�{P uiH�{@ �����1�A�   �D$k���$�   H���[���H�L$PD���    L�	A�Q��A�������H��$�   �m �����f��$�   ����L��H���Q���������  H�{@ �y���H�{P �n����r���H��PP�����H��PP�����H;|$H�����H��$�   H�x���   �|$k �7  H��$�   H�x� t>�D$l@��E��H��$�   H��E����  H�SI��H�K�� ��uH��$(  �E��uzH�T$8H��$0  虴  L�d$pH��$�   �9���H��PH�����H��PH����H��PH�����L;l$`�L���M�������H��$   �@�D$`%   A��@�������9sX������x���H�|$8E1��0   H���A��H�������H��$�   H���A�    H��L�B�I�P�HD�L9�LF�1���  �������$�   H���q���H�S8f9�����H�C@H��$�   H�D$H�.k A�����A�   fD��$�   �I�����$�   H���$���H�SHf9����H�CPH��$�   H�D$H��j A�����A�   �D$kfD��$�   �����f�E�������H��$�   H�x����������H��PHD��� ����|$j@���l�����$�   �^�����$�   ������K���H��PH����H��$�   �P���ye�80������@���yIH�L$8A�   E1�1��D$ -   �
�  H��$�   �@������y���E1����u      ��A�������E�������H�L$8��  �H�L$8���  H��$�   �E1�����H��$�   H��H��$�   H��H�H���  H��$�   H��H�H���  H���+���H��$�   H���א�������������SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����SH��`�Ao�AoH�)D$@L�L$@H��H��$�   )L$PL�D$PH�L$8H��$�   H�L$0H��$�   H�L$(��$�   �L$ H���PH��H��`[Ð����AVAUATUWVSH��   )�$�   )�$�   H��$  D��$  �Ao �Ao9H��I��)D$@H��$(  H���   � H��$�   1�1�I��I���o�  H�L$pE��H��$�   ��   H��$�   foL$@H�t$ L��H�D$0H��$   L�L$PL�D$`)L$`)|$PH�D$(����H�L$xH�D$pH�L$xH��$�   H�D$pH�D$@fot$@f�t$xH�q�H��t=E1�H��H���s6  H��@�����   H��$�   L��I�$L�L�2�PXH��$�   3�������A���~s(�$�   H��(�$�   H�İ   [^_]A\A]A^�H��$�   foT$@H�t$ L��H�D$0H��$   L�L$PL�D$`)T$`)|$PH�D$(����������     H��H���$�  �|���H���G$  �=���H��H��$�   H��H�H���  H���3������ATUWVSH��   )�$�   D��$�   �Ao �Ao9H��$   H��$�   H��H��)D$@1�1�I��蒨  H�L$pE��H��$�   ��   H��$�   foL$@H�|$(H��H�D$0H��$�   Lv      �L$PL�D$`)L$`)|$PH�D$ �;���H�D$pH�T$xH�D$@fo|$@H�T$xf�|$xH�D$p�0� H��$�   I��I��H��$�   H��$  �m� H��$�   >�������A���~d(�$�   H��H�Ġ   [^_]A\�H��$�   foT$@H�|$(H��H�D$0H��$�   L�L$PL�D$`)T$`)|$PH�D$ �:����:���D  H��H���t�  �H��H��$�   H��H�H��k�  H���������SH��P�Ao H�H��)D$@E��H��$�   L�D$@H�L$0��$�   �L$(H��$�   H�L$ H���PH��H��P[Ð������������SH��`H��$�   �Ao �(H��)D$PE��H�L$@H�H�L$0��$�   L�D$P�|$@�L$(H��$�   H�L$ H���PH��H��`[Ð�SH��@�D$x�Ao�D$ L�D$0H��E��H��$�   )L$0L�L$pH�L$(H��t�1	  H��H��@[��     �[  H��H��@[Ð�UAWAVAUATWVSH��   H��$�   )}���   �Ao8�E�H���   H��H�MpH��H�UxD�M��(H���   �}�H���   �� H���j H��@I��H�\$0I����� �m�A�@   H��H�E�D$     H�u�}�L�e�H��L��� L�d$(�_� ��?~O�XHc�H��H�������H)�L�|$0M���g� �m�L�d$(A��L���D$     H��L�W� H�E�}��� Hc�E1�H��L�}�H��M����  L�eA�D$�����   A�E8<t ����   I�E H�����H�@8H9���   I��L��L�������E�)}�L�EЀ}� H�t$(L���   H�Ux�D$ H�MptA�|  H�M�������A���~ZH���� H�Ep(}H�e([^_A\Aw      ]A^A_]�f�     �{   �f�     H����  L�e�=���L���'����A���f�H��L���$�  �f�M��L��L��M����A���H���H��H�EL��H�H���  H����� H���$�������AWAVAUATUWVSH��   I� I�xH�D$8��$   M���   L��H��$   L����D$T�D$P�6 H��_ I�������I��H���   H�@N�$�I�$H����  H��$(  L�(�CdA8E M�e��k  �C\��$�   H�C8H�D$`H�C@H�D$@M�M9�v.I�O0L��A�U �Qu� ��QtGH��I9�u�M)�uAH��$   H�F    @��H�t$8H�xH�0H�ĸ   [^_]A\A]A^A_�fD  I��M)�t�H��$�   1�1�L��$�   I��H�D$H臢  K�$L��L�t$XH��$�   �N�  �CXE��A)�E����   ��EH�H�{ �   G�?1�L��L�t$XH��$�   Mc�L�@��D$     ���  Ic�H��$�   L�D�s"H�D$hH�CH�D$pH�CH�D$x�A����  H�D$hD��L�l$ L�L$pL�D$xH�D$(�+� H��$�   I�ƋA�����  L�I�L��H)�M��I)�L9���  H�L$XE1��_�  �CX���t  �FH��$�   L�t$@����   Lr����L$p�  L��$�   1�1��J�  H�L$HK�6H��$�   ��  H�NL��$�   �|$pM�|$L�-3| H�L$h��L9���L)�!��D$PI�ΈT$x�D$PA�<$��   A�$IcD� L���f.�     �C`M�䉄$�   �����H�CHI��H�D$`H�CPH�D$@����f�H�|$@ txH�D$`H�L$H�趷  �d@ �FtZH�S(L�C0H�L$H�(�  x      �FfD  �|$x �v  D�D$PL��H�L$H�C�  �!��|$x t���    H�T$XH�L$H�Ѩ  �I��M9�����H�D$@H����   H��$�   H�\$hH�B�H9�wq@��Hc�uH�L$8I��H��P`H��$�   H9�@��H�\$8H�J�1�@��@��H��$�   ��H��$�   H��$�   H��趣  H��$�   H��H�H�袣  ����H)Ã|$p D�D$TI���P  H�L$HD�D$ 1�E1���  H��$�   H�D$h�R���Ls0������    H�T$`L�@�H�L$HH���٦  ����@ L�t$X�S!L���/�  E����   LcCXIc�L��L�褦  �[����T$PH�L$H��  �����p   ��* H���@    L��H��> H�C    H��H�1�H�C    f�C �C" H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co �F� H���   H��M���� I�$�����H�L$XMc�L���+�  ����H�L$HH���	�  ����A��D�CeIc�L�|$XL����  M��L��L��螥  �U���H�L$X蟝  H��$�   �����H�L$X舝  H��$�   �����H�tx I��H�Rx �5� H��$�   H��H��$�   H��H�H�薡  H��$�   H��H�H�股  H������H��$�   H����H���e+ H�H���P�2 H���O+ ��H���e- H���m����������������AWAVAUATUWVSH��   I� I�xH�D$8��$   M���   L��H��$   L����D$T�D$P�v� H�Y I���7���I��H���   H�@N�$�I�$H����  H��$(  L�(�CdA8E M�e��k  �C\��$�   Hy      �C8H�D$`H�C@H�D$@M�M9�v.I�O0L��A�U �Qu� ��QtGH��I9�u�M)�uAH��$   H�F    @��H�t$8H�xH�0H�ĸ   [^_]A\A]A^A_�fD  I��M)�t�H��$�   1�1�L��$�   I��H�D$H�Ǜ  K�$L��L�t$XH��$�   莰  �CXE��A)�E����   ��EH�H�{ �   G�?1�L��L�t$XH��$�   Mc�L�@��D$     ��  Ic�H��$�   L�D�s"H�D$hH�CH�D$pH�CH�D$x�A����  H�D$hD��L�l$ L�L$pL�D$xH�D$(�k� H��$�   I�ƋA�����  L�I�L��H)�M��I)�L9���  H�L$XE1�蟰  �CX���t  �FH��$�   L�t$@����   Lr����L$p�  L��$�   1�1�芚  H�L$HK�6H��$�   �T�  H�NL��$�   �|$pM�|$L�-_u H�L$h��L9���L)�!��D$PI�ΈT$x�D$PA�<$��   A�$IcD� L���f.�     �C`M�䉄$�   �����H�CHI��H�D$`H�CPH�D$@����f�H�|$@ txH�D$`H�L$H����  �d@ �FtZH�S(L�C0H�L$H�h�  �FfD  �|$x �v  D�D$PL��H�L$H胣  �!��|$x t���    H�T$XH�L$H��  �I��M9�����H�D$@H����   H��$�   H�\$hH�B�H9�wq@��Hc�uH�L$8I��H��P`H��$�   H9�@��H�\$8H�J�1�@��@��H��$�   ��H��$�   H��$�   H�����  H��$�   H��H�H���  ����H)Ã|$p D�D$TI���P  H�L$HD�D$ 1�E1��2�  H��$�   H�D$h�R���Ls0����z      ��    H�T$`L�@�H�L$HH����  ����@ L�t$X�S!L���o�  E����   LcCXIc�L��L���  �[����T$PH�L$H�A�  �����p   �"$ H���@    L��H�.8 H�C    H��H�1�H�C    f�C �C" H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Co �V� H���   H��M���T� I�$�����H�L$XMc�L���k�  ����H�L$HH���I�  ����A��D�CeIc�L�|$XL���,�  M��L��L���ޞ  �U���H�L$X�ߖ  H��$�   �����H�L$X�Ȗ  H��$�   �����H��q I��H��q �u� H��$�   H��H��$�   H��H�H��֚  H��$�   H��H�H��  H�������H��$�   H����H���$ H�H���P�G+ H���$ ��H���& H�������������������SH��P�Ao H�H��)D$@E��H��$�   L�D$@H�L$0��$�   �L$(H��$�   H�L$ H���PH��H��P[Ð������������SH��`H��$�   �Ao �(H��)D$PE��H�L$@H�H�L$0��$�   L�D$P�|$@�L$(H��$�   H�L$ H���PH��H��`[Ð�SH��@�D$x�Ao�D$ L�D$0H��E��H��$�   )L$0L�L$pH�L$(H��t�	  H��H��@[��     �  H��H��@[Ð�UAWAVAUATWVSH��   H��$�   )}���   �Ao8�E�H���   I��H��H�UxH��D�M��(H���   �}�H���   �#� H����� H��@I��H�\$0I����� �m�A�@   H��H�E�D$     H�u�}�L�m�H��L�Js L�l$(�p� {      ��?~R���E�H�H��H��������H)�H�\$0I���v� D�E�L�l$(H��H���m��D$     H�EL��r �}��� Hc�E1�H��L�m�H��M���+  L�MA�A�����   I�M�L��L���PX�E�)}�L�E�L���}� H�t$(L���   H�Ux�D$ t8�s  H�M�������A���~BH����� �(}L��H�e([^_A\A]A^A_]��[   ��f�     H���  L�M�n���H��L���c  �H���H��H�EL��H�H��Y  H���a� H���������������AWAVAUATUWVSH��   I� I�xH�D$8��$   M���   L��H��$   L�����D$xf�D$T��� H�NO I���V���I��H���   H�@N�,�I�] H����  H��$(  �KdL�(fA9M I�E�t}�S\��$�   H�S8H�T$XH�S@H�T$@M�$L��M��   M�LE A�R(L)�I��I��I��ukH��$   H�F    @��H�t$8H�xH�0H�ĸ   [^_]A\A]A^A_��     �S`H����$�   H�SHH�T$XH�SPH�T$@I�ULE��s���@ H��$�   1�1�I��H�D$H�G  L��H��$�   H��$�   H��H�D$`�#  �CXE��A)�E����   ��EH�H�{ �  H��$�   G�$61�H�L$`Mc�M��L�@��D$     ��  H�SM�H��$�   H�T$hH�SH�T$p�S$�T$|�A����  L�L$hL�d$(L�D$pL�l$ �T$|��� H��$�   I�ċA����  L�I�L��H)�H��M��I)�L9��  H�L$`E1���#  �CX���c  �FL�t$@��   �T$pH��$�   Lr����
  L��$�   1�1��	  H�L$HK�6H��$�   |      �"  H�NL��$�   �|$pM�|$L�-o H�L$h��L9���L)�!��D$TI�ΈT$|�D$TA�<$��   A�$IcD� L���f�     H�|$@ txH�D$XH�L$H��F$  �d@ �FtZH�S(L�C0H�L$H��  �FfD  �|$| ��  D�D$TL��H�L$H�  �!��|$| t���    H�T$`H�L$H�  �I��M9��P���H�D$@H����   H��$�   H�\$hH�B�H9���   @��Hc�uH�L$8I��H��P`H��$�   H9�@��H�\$8H�J�1�@��@��H��$�   ��H��$�   H��$�   H���"  H��$�   �������A��������H��H����  �����    H)Ã|$p D�D$xI���i  H�L$HD�D$ 1�E1��5  H��$�   H�D$h�9��� Ls0������    H�T$XL�@�H�L$HH���i  �����@ L�d$`�S"L���"  E���  LcCXMc�L��K�Tu �2  �j����T$TH�L$H�o"  ����f.�     ��   �6 H���@    L��H�b. H�C    H��H�H�C    �C  �C"    H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz �9� H���   H��M���g� I�] �����H�L$`Mc�L����  ����f�     H�L$HH���  ����A��D�CfIc�L�t$`L���v  M��L��L���  �P��� H�L$`�V  H��$�   �����f�     H�L$`�6  H��$�   �����H�Bk I��H� k �s� H��$�   H��H��$�   H��H�H���  H��$�   H��H�H��  H�������H��$�   }      H����H��� H�H���P�E! H��� ��H��� H�����������������AWAVAUATUWVSH��   I� I�xH�D$8��$   M���   L��H��$   L�����D$xf�D$T�� H�~H I���v���I��H���   H�@N�,�I�] H����  H��$(  �KdL�(fA9M I�E�t}�S\��$�   H�S8H�T$XH�S@H�T$@M�$L��M��   M�LE A�R(L)�I��I��I��ukH��$   H�F    @��H�t$8H�xH�0H�ĸ   [^_]A\A]A^A_��     �S`H����$�   H�SHH�T$XH�SPH�T$@I�ULE��s���@ H��$�   1�1�I��H�D$H�g  L��H��$�   H��$�   H��H�D$`��  �CXE��A)�E����   ��EH�H�{ �  H��$�   G�$61�H�L$`Mc�M��L�@��D$     �
	  H�SM�H��$�   H�T$hH�SH�T$p�S$�T$|�A����  L�L$hL�d$(L�D$pL�l$ �T$|�� H��$�   I�ċA����  L�I�L��H)�H��M��I)�L9��  H�L$`E1���  �CX���c  �FL�t$@��   �T$pH��$�   Lr����
  L��$�   1�1��)  H�L$HK�6H��$�   �  H�NL��$�   �|$pM�|$L�-h H�L$h��L9���L)�!��D$TI�ΈT$|�D$TA�<$��   A�$IcD� L���f�     H�|$@ txH�D$XH�L$H��f  �d@ �FtZH�S(L�C0H�L$H��  �FfD  �|$| ��  D�D$TL��H�L$H�#  �!��|$| t���    H�T$`H�L$H�  �I��M9��P���H�D$@H����   H��$�   H�\$~      hH�B�H9���   @��Hc�uH�L$8I��H��P`H��$�   H9�@��H�\$8H�J�1�@��@��H��$�   ��H��$�   H��$�   H���B  H��$�   �������A��������H��H���  �����    H)Ã|$p D�D$xI���i  H�L$HD�D$ 1�E1��U  H��$�   H�D$h�9��� Ls0������    H�T$XL�@�H�L$HH���  �����@ L�d$`�S"L���  E���  LcCXMc�L��K�Tu �R  �j����T$TH�L$H�  ����f.�     ��   �V H���@    L��H��' H�C    H��H�H�C    �C  �C"    H�C(    H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    �C`    �Cz 詔 H���   H��M��臲 I�] �����H�L$`Mc�L����  ����f�     H�L$HH���  ����A��D�CfIc�L�t$`L���  M��L��L���8
  �P��� H�L$`�v  H��$�   �����f�     H�L$`�V  H��$�   �����H�bd I��H�@d �� H��$�   H��H��$�   H��H�H���  H��$�   H��H�H���  H������H��$�   H����H���� H�H���P�e H��� ��H���� H�������������������+   �����������1�Ð������������1�Ð������������H��(�   H9�t$H�I1��9*tH�R1��:*��H���������H��(Ð������������H)�H������@H��   �M�ÐH�Ð�����������H�Ð�����������SH�� H��@�H�˅�~E1�E1�1��  H      ��@�����H�� [ÐWVSH�� H�ˉ׉�1���  H��H��H�@t1�H��t7�    f�tQH��H9�u�1��A    H�f�TYH�� [^_�f�     f�y�ؐ���������UWVSH��(H��H��1�H)�H��H��H���O  H��L�HH��t5H��u1��C    H�;f�D3L��H��([^_]�L��I��H�����I�����E f�C�Ɛ��UWVSH��(H��H��tH��thH��1�H)�H��H��H����  H��L�HH��t;H��u#1��F    H�>f�DL��H��([^_]�fD  L��I��H���~��I�����E f�F��H��V 臾 �������UWVSH��(H��H��tH��thH��1�H)�H��H��H���E  H��L�HH��t;H��u#1��F    H�>f�DL��H��([^_]�fD  L��I��H���~��I�����E f�F��H�V ��� �������H�i> Ð�������I)�L��H��H��tH��u��}��fD  �f�Ð��������I)�L��H��H��tH��u��}��fD  �f�Ð��������I)�L��H��H��tH��u��V}��fD  �f�Ð��������I)�L��H��H��tH��u��&}��fD  �f�Ð��������H��(H�H�P�H9P�rH��(�f.�     1��  �H��(�H��� �H��(�� �ATUWVSH�� H��l$pI��H��L��H����������L�H+P�I9�wOL���6  H��tH�1�H��J�`t"f�f�<PH��H9�u�H��H�� [^_]A\�D  f�(H��H�� [^_]A\�H��S �c� ���UWVSH��(H�\$pL��I��H��H����  H��tH�H��H�xt L�H���|��H��H��([^_]À      �     �E f�H��H��([^_]Ð���������������������������VSH��(H�L�@�H��H��L9�s�P���x����H�H�XH��([^�H�R ��� ��SH�� H��P�H�˅�x�Y���H�H�P�H�PH�� [Ð��������� ������������������A��~Ð� �������������AH�AÐ�����H�AÐ����������H��; Ð��������A����Ð��������A    Ð�������1��A    H�f�DQÐ�������������D�AH�AE��x�� H�A�f.�     E1��   ��������VSH��(H��H�	L�I��H�V�e   1�H��H�L�KH��t L� H��t:H�VL���>z��I��H�H� H�1��C    f�DL��H��([^�f�     �Vf�S�   �͐SH�� H��������H9�H��weH9�vEH�H9�HB�H�LL�A I��   v-H9�s(A���  �   L)�H��H�H9�HG�H�L�H�L	�e
 H�X�@    H�� [�H��P 蘺 ��������VSH��(H�H��H�H�P�H�Y���xH���=���H�H�XH��([^Ð��������������VSH��(H��H�
H�֋A���xH������H�H��H�H��([^Ð�H�D�@�E��y�@�    L�E�H�E��yA�@�    L�H�Ð�SH�� H��P�H�˅�x����H�H�� [�E1�1�H�L�@��?  ���������������VSH��(E1�A�   H��H+H��H��H���  H��@�����H�H��([^Ð��������VSH��(I)�H��H��I��uH��([^�D  H+E1�H��H��H���  H�H��B�����H��([^Ð�������      SH�� H�L�H�H��L��H)�L9�LF�L9�wE1�H���t  H��H�� [�H��N I��H�7O �� �����SH�� H��P�H�˅�x����H�H�� [�VSH��(H��H��H���v��H��H��I��H��([^�   ��������UWVSH��(M��H��H��L��txH��������H�H�X�H)�I9���   L�H;X���   H9�wH�P�H�PH9�vNH��H���  H�H�P�H��H�PtTL�?H����v��H�1��@�    H�X�f�XH��H��([^_]�fD  H��H��H)��b  H�H�P�H�H��H�Pu��U f��D  �@���H��b����H�gN 蔷 ����UWVSH��(H�H�p�H��H��H��tLH�H�h�H�H;h�vHH��H����  H�H��H�H�H�H�Ht7L�6�v��H�1��@�    H�h�f�hH��H��([^_]Ë@�����D  �f��͐�������UWVSH��(H�H�X�H��H��I9���   L)�L9�IG�H��taH�H�h�H�H9h�r�@���~H��H��L�D$`�<  L�D$`H�H��J�@H�H�H�H�Ht/L��fu��H�1��@�    H�h�f�hH��H��([^_]�fD  �f���H�M I��H��K �r� ��H��H�L�@�����SH�� H��H��t	E���
   H��H�� [ÐATUWVSH�� H��������H��H�H��E��D��H�r�H)�H9�rwH�H;r�vXH��H���]  H�M H��H�A�H�AtKH��t1�@ f�<BH��H9�u�1��A�    H�q�f�qH�� [^_]A\��    �B������    fD�"��H�1L �^� ��������������H��(�'���H��H��(Ð��������������VSH��(H��      �H��H���4s��H��H��I��H��([^�   ��������VSH��8H�L��I��H��L�@�H��������H9���   L9�vH�t$ 1�H���c���H��8[^�J�@I9�w�@���~H�L�@��� H�	L�6L��H)�H��H9�v;H��tH��tPH��tL���Ks��H�1��A�    H�q�f�qH���f.�     H��tH��t�L���s��H����     A�f��H��J �� �����������VSH��8H�2H91H��t'�V�H�N�H�A��x"�� H��������A���~H�3H��H��8[^�H�T$/E1��!���H����H���# �֐H��(L�I�R�H��L)�L9�IG�I9�wK�BI��H��(����H�I I��H�+J 蝹 �������������H��H�L�@�Q����H��8H�H�@�E��I��1�D�D$ I���?���H��8Ð���������H+M�HM� H���   ��������������VSH��8A�   H��H+E��H��D�D$ E1�H��H�������H��@�����H�H��8[^�H��8H+E��H��D�L$ M��E1������H��8Ð�����������WVSH�� H��L��H��L���p��I��H��H��I��H�� [^_�    ATUWVSH��0H��H�L��H��L�J�L9��V  H��������L)�H9��4  L9�v"M��H�l$ E1�H��H������H��0[^_]A\ÐJ�JI9�wՋB����H��L��I��H+1E1�H��Y  L�L�d- I�1I�J�"L9�w#H����   H���~   M��L���p��H���L9�r%H���   H��tZM��H��L���\p��H���h���H)�H��H��H��tLH��tL��I���5p��I��K�!H)�I�9H��t@H��tL�D- �p��f��      H�������fA�H�������fA��� fA�H��������f�H�������H�zG �� H�nG I��H�vF �� �M� M�H��d�������H��(M�L�T$PM�C�L��M��I)�M9�MG�L9�wM�CH��(�.���H�G M��I��H�F 襶 �����H��8H�H�@�E��H9�wD�L$ M��E1��\���H��8�H��E I��I��H��F �^� ��������������VSH��(H��H�
H�֋A���xH�������H�H�A�H�AH�H��H��([^Ð���������E1��   ��������H��(I��������H�L9�H�@�w8H9�w#rH��(�f.�     H)�E1�I��H��(�  H)�E��H��(�n���H�ZF �r� ��I��tM��u�@ M��8n���     �f�Ð��������H��H�Ð��������H��@���y�D  ����������������I��tM��u�@ M���m���     �f�Ð��������H�D$(I)�H+L)�H��I��H�D$(H����  ���������������UWVSH��8H��H��L��L��L��H)��l��H+I��I��H�D$ I��H��H��H���  H��8[^_]Ð��������H�D$(I)�H+L)�H��I��H�D$(H���O  ���������������I)�H+I��H���/  ���������������H��8M�	I)�I�A�H+I��H�D$ H����   H��8Ð���������H�D$(I)�H+L)�H��I��H�D$(H����   ���������������H�D$(I)�H+L)�H��I��H�D$(H���   ���������������H��8I�AH�I)�H+H��H�D$ M�	I��H���i   H��8Ð����D$(I)�H+�D$(I��H���F�      ��������UWVSH��8H��L��H��L��L���,k��I��I��H��H�D$ H���   H��8[^_]Ð����AVAUATUWVSH��@H��$�   H��L��H��H�L�H�L9��<  L��H)�H��������L9�IG�L)�H�H9��,  H9�v+I��H�l$ H��I��H��� ���H��H��H��@[^_]A\A]A^�J�HH9�w̋@����H�L�l- L�4?J�)N�0L9���   L�N�@L9�rAH)�H��L�$)I)�H��H��I��I���  H�J�aL�H��tsH��t�M����j���t����L�l$?E1�M�������H�l$ I��H��I��H��I���g���H�Ƹ�����A�D$����3���I�L$��� �$����H)�H��I���n���f��f�����H�A I��H�B 蟱 H�B �c� I�L$�H��L�������H���+��������������H��8M�	I�A�H�D$ �;���H��8Ð�����SH�� I�L�T$PL�\$XL�K�L��L)�L9�IG�M9�wN�SH�D$PH�� [�����H��A M��H�t@ ��� ���������������H��(H�D�\$PL�P�L��H)�L9�LF�L9�wD�\$PH��(����H�(@ I��M��H�A 覰 ������SH��@H��H�	H;Q�tTH�A�H9�HB�H��I��H�T$?I)�����H��������Q���~H�H��@[�fD  H��H�D$(�� H�D$(�܋A���~�H�렐��������������H��(E1�H�H�@�H�P�H9�wA�   H��(�J   H� @ I���H�X? �� ���H��E��tH��t1�fD�AH��H9�u�ÐfD�Ð����������AWAVAUATUWVSH��8H�I��H�P�L��H��O�, L)�L��H�L)�I��H�P�H9�w�@���      ���   H�H�P�L�D$/H������M��I��uaH�pH�M��t"J�hL�I��I�Lo��   O�6��g��H��������P���~rH�71��F�    H�^�f�^H��8[^_]A\A]A^A_�H�I�wI��tOO�$H��H���g��H��M��H�1t�M9�t�J�nL�I��H�nt=O�6�Lg��H�7�H�H���� �@ �fA�W�=��� �f��V���D  �f��W��������WVSH�� H�H��H�H��H�YH;X�w�@���~H��H������H�H�P�f�<P1��@�    H�X�f�XH�� [^_Ð������������SH��0H�L�D$/H��H�1�1�����1��@    H��H�@�    f�H�H��0[Ð��VSH��(H��H��H������H��tH��L�D$P�e��L�D$PH�CE1�H���7���H�H��([^Ð������������SH�� L��H��E1�H��J�BI������H�H�� [Ð���������SH�� H��I��1�1������1��@    H��H�@�    f�H�H�� [Ð����������SH��0H�D�@�H��H�H�H�QE��x��H�H��0[��    H�T$/E1������H�H��0[Ð���������SH�� H�M��L�H�H��J�HM9�wJ�@E1�M�������H�H�� [�H�h= H��; �j� ����������SH��0H��H�
L�Q�L��L)�L9�IG�L�M9�H�AwJ�AE1�L�D$/�g���H�H��0[�H�	= M��H�}; �� ��������SH�� H��H�
L�Q�L��L)�L9�IG�L�M9�H�AwJ�AL�D$PE1�����H�H�� [�H��< M��H�; 訫 ��������SH�� E1�H�BH��H�
H�A�5���H�H�� [Ð����      ��������SH��01�L�D$/H��1��
���1��@    H��H�@�    f�H�H��0[Ð��������SH�� H��H��A��M�������H�H�� [�SH�� H��H��L��M��E1��7���H�H�� [Ð�������������SH�� H��H��L��M��E1��w���H�H�� [Ð�������������SH�� H��H��L��M��E1������H�H�� [Ð�������������SH��0H�L�D$/H��H�1�1�����1��@    H��H�@�    f�H�H��0[Ð��VSH��(H��H��H������H��tH��L�D$P�b��L�D$PH�CE1�H������H�H��([^Ð������������SH�� L��H��E1�H��J�BI������H�H�� [Ð���������SH�� H��I��1�1��\���1��@    H��H�@�    f�H�H�� [Ð����������SH��0H�D�@�H��H�H�H�QE��x��H�H��0[��    H�T$/E1��s���H�H��0[Ð���������SH�� H�M��L�H�H��J�HM9�wJ�@E1�M���F���H�H�� [�H��9 H�_8 �� ����������SH��0H��H�
L�Q�L��L)�L9�IG�L�M9�H�AwJ�AE1�L�D$/�����H�H��0[�H��9 M��H��7 舨 ��������SH�� H��H�
L�Q�L��L)�L9�IG�L�M9�H�AwJ�AL�D$PE1�����H�H�� [�H�)9 M��H��7 �(� ��������SH�� E1�H�BH��H�
H�A����H�H�� [Ð�����������SH��01�L�D$/H��1�����1��@    H��H�@�    f�H�H��0[Ð��������SH�� H��H��A��M���i���H�H�� [�SH�� H��H��L��M��      �E1�����H�H�� [Ð�������������SH�� H��H��L��M��E1������H�H�� [Ð�������������SH�� H��H��L��M��E1��W���H�H�� [Ð������������������H�	��A���~�H���%� ����������H�	��A���~�H���� �����H��(�g���H��H��(Ð��������������VSH��(H��H��H���t^��H��H��I��H��([^�H������������+��������������SH�� H��H�H��L�@����H��H�� [�SH��0A�   H�L�@���H�ˉT$ 1������H��H��0[Ð���VSH��(H�H�֋P�H�˅�x����H�H�pH��([^Ð������VSH��(H��H��H���]��H��H��I��H��([^����������������������������H��H�L�@������WVSH�� H�H��H�H��H�YH;X�w�@���~H��H�������H�H�B�f�<B1��B�    H�Z�f�ZH��H�� [^_Ð���������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���Z H���   H����r H���   H����r H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�W���   H�EH�UH�GH��([^_]Ð�����������UWVSH��(H�iH��H��H����c 1�H��Hǃ�       f���   H�� H�H��(H�CH�GHǃ       Hǃ      Hǃ      H�CH�Hǃ      H�p�H�H���W H���   H���q H���   Hǆ�       H���   ���   ���   ���   Hǃ       ���   H��� H�G    H��      H��PH�CH��(H�CH��([^_]�H��H��� H��H�PH�S�c H��������������������UWVSH��(H�-	� H�qH��H��H���b 1�H�+H��f���   H�E(H��Hǃ�       Hǃ       Hǃ      Hǃ      Hǃ      H�CH�C    ��q H�� H��H��H�CH��(H�C��q H��� H�H��PH�CH��(H�CH��([^_]�H��H��� H��H��H�C�b H������H�+H��H�C    �ѐ�������������WVSH�� H�=
� H�qH��H���a 1�H�;1�f���   H�G(H��Hǃ�       Hǃ       Hǃ      Hǃ      Hǃ      H�CH�C    ��p H�� 1�H��H�CH��(H�C��p H��� H�H��PH�CH��(H�CH�� [^_�H��H�� H��H��H�C�a H������H�;H��H�C    �ѐ����ATUWVSH�� H�BH��H��H�H�JH�P�M��H�I�PH�SH�x�I� H�H�h�H��L�H����T H���   H����n H���   Hǅ�       H���   ���   ���   ���   HǇ�       ���   H�FI�D$    H�CH�@�H�V H�TH�H�H�@�H�V(H�H�F0H�CH�� [^_]A\Ð�����WVSH�� H�BH��H�H��H�JH�P�L��H�L��H�C    H�H�H��Vo H�FH��H�CH�@�H�LH�F H��6o H�H�H�@�H�V(H�H�F0H�CH�� [^_�H�VH�H�R�H�NH�H��H�C    聰���VSH��(H�BH��H�H��H�JH�P�H�1�H�C    H�H�H��n H�F1�H�CH�      �@�H�LH�F H��n H�H�H�@�H�V(H�H�F0H�CH��([^�H�VH�H�R�H�NH�H��H�C    ������������SH�� H�L� H�AH�� H��H�H�,} H�IH�A�    H��H��$_ H��H�� [�'� �������H�� H�AH��� H��H�A�H��| H�A�    H��H���^ �����������H�H�H�@�L�B(L�H�B0H�AH�BH�AH�@�L�B L�DH�BH�H�@�H�RH�H�A    Ð����UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���#S H���   H����k H���   H����k H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�U���   H�GH�WH�EH��H��([^_]Ð��������VSH��   E1�H��H��H�L${H���a$  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R`�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q �m H��H�Ĉ   [^�蜑 H��H��t �.� H�H�p�HރN �Fu7�5� ��� H�HX�K �Cu�� �� H���� H�������� H����� H���������������������VSH��   E1�H��H��H�L${H���#  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R�T$|��uH��H�Ċ      �   [^ÐH�H�H�H�Q �nl H��H�Ĉ   [^��L� H��H��t ��� H�H�p�HރN �Fu7��� ��� H�HX�K �Cu�X� �S� H���� H���ë���>� H���� H��讫����������������VSH��   E1�H��H��H�L${H����!  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�RP�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q �k H��H�Ĉ   [^���� H��H��t �� H�H�p�HރN �Fu7�� ��n� H�HX�K �Cu�� �� H���k� H���s������ H���V� H���^�����������������VSH��   E1�H��H��H�L${H���q   �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�RX�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q ��i H��H�Ĉ   [^�謍 H��H��t �>� H�H�p�HރN �Fu7�E� ��� H�HX�K �Cu�� �� H���� H���#����� H���� H��������������������VSH��   E1�H��H��H�L${H���!  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�RH�T$|��uH��H�Ĉ   [^Ð�      H�H�H�H�Q �~h H��H�Ĉ   [^��\� H��H��t ��� H�H�p�HރN �Fu7��� ���� H�HX�K �Cu�h� �c� H����� H���ӧ���N� H���� H��辧����������������VSH��   E1�H��H��H�L${H����  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R(�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q �.g H��H�Ĉ   [^��� H��H��t �� H�H�p�HރN �Fu7�� ��~� H�HX�K �Cu�� �� H���{� H��胦����� H���f� H���n�����������������VSH��   E1�H��H��H�L${H���  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q ��e H��H�Ĉ   [^�載 H��H��t �N� H�H�p�HރN �Fu7�U� ��.� H�HX�K �Cu��� ��� H���+� H���3����� H���� H��������������������VSH��   E1�H��H��H�L${H���1  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R0�T$|��uH��H�Ĉ   [^ÐH�H�H�H�      �Q �d H��H�Ĉ   [^��l� H��H��t ��� H�H�p�HރN �Fu7�� ���� H�HX�K �Cu�x� �s� H����� H�������^� H����� H���Σ����������������VSH��   E1�H��H��H�L${H����  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R �T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q �>c H��H�Ĉ   [^��� H��H��t �� H�H�p�HރN �Fu7�� ��� H�HX�K �Cu�(� �#� H���� H��蓢���� H���v� H���~�����������������VSH��   E1�H��H��H�L${H���  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R8�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q ��a H��H�Ĉ   [^��̅ H��H��t �^� H�H�p�HރN �Fu7�e� ��>� H�HX�K �Cu��� ��� H���;� H���C����� H���&� H���.�����������������VSH��   E1�H��H��H�L${H���A  �|${ t|H��D$|    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$(L�D$PH�D$@    L�L$PL�L$@H�t$0H�D$ A�R@�T$|��uH��H�Ĉ   [^ÐH�H�H�H�Q �`�       H��H�Ĉ   [^��|� H��H��t �� H�H�p�HރN �Fu7�� ���� H�HX�K �Cu�� �� H����� H�������n� H����� H���ޟ����������������WVSH��0H�H�@�H��H��H���   H��t_�{8 tD�KCH��H��H��0[^_�R   f�H��L�D$(�3<��H�A�
   H�c>��L�D$(H�@0H9�t��
   H����L�D$(D����{� �����������ATUWVSH��0H��H�A    H��M��H�L$/A�   H��D���O  �|$/ u8M���?  � H�{ u�   H�H�H�H�Q �_ H��H��0[^_]A\�H�@��H�@�H���   H�FH9FwQ H�H���PHH�SH�JL9�|Hf.�     ����  M����   � H�{ u��z���H��H�FH9�s�H�S� H�JL9�}��t39���   H���G�H�FH�VH�CH9�r�H�H���PP�����   �   M��~� H�{ uf������H��H����   �� H�H�p�HރN �F��   �� M�������fD  H�SH�������H��H��0[^_]A\�D  �������H��H��0[^_]A\�f.�     1��d���M��~!� H�{ t�   �p���H�FH�V�����H��u�   �T����� H�HX�K �Ct�� �� H���� H�������� H����� H����������������������WVSH�� H�H�@�H��H��H���   H��tP�{8 tD�CCH��H��H�� [^_�B   f�H���X9��H�H��;��A�
   H�@0H9�t˺
   H����D���誀 ����������UWVSH��8�      H��H�A    H��D��H�L$/A�   H���  �|$/ t`H�@��H�@�H���   H�FH9Fvp� ��9�t:H�C(H;C0s}�H�C(H�FH�VH�GH9�sxH��H�FH9�v7���9�u�H� u�   H�H�H�H�Q ��[ H��H��8[^_]� H�H���PH�����u�H�҃����H�H���Ph����x����H�H���PP���t�H�FH�V�u���H��H��u�#� H�Hx�O �Gt#�� �� H�H�H�H��I �At�� �� H���� H���
������ H� �$����6���H����� H�����������VSH��8A�   H��H�A    H��H�L$/H����  �|$/ u2H�{ u�   H�H�H�H�Q ��Z H��H��8[^�f.�     H�H�@�H���   H�AH9Av'�H��H�AH�C   �H�{ t�H��H��8[^ÐH��PP���uH�{҃���뀉���H��H��u��� H�HX�K �Ct#�~� ��� H�H�p�HރN �Ft�`� �[� H����� H���˙���� H�{ �����"���H���� H��覙��������SH��0A�   H��H�A    H�L$/H���  �|$/ ��   H�H�@�H���   H�QH9Qv�H��H�QH�C   H��0[�H��PP���u�H�{҃���H�HX�S H���VY �����H��0[�H��H��t0��� H�H�P�HڃJ �BuG��� @ H�{ uú   ��� H�HX�K �Ct�7� �2� H���� H��袘���� H���� H��荘���������������SH��@A�   H��HǏ      A    H�L$?H���  �|$? tvH�H�@�H���   H�AH9Av� H��@[�@ H��PH���u�H��D$,HZ�S H�ك��LX �D$,��H��H��t$��� H�HX�K �Cu>��� f��������� H�HX�K �Ct�>� �9� H���� H��詗���$� H���� H��蔗������WVSH��0H��H�A    H��L��H�L$/A�   H���  �|$/ t$H�I��H��H�@�H���   H��P@H9�H�CuH��H��0[^_�H�H�H�HًQ ���ZW H��H��0[^_�H��H��t ��� H�H�x�H߃O �Gu7��� ��� H�HX�K �Cu�K� �F� H���� H��趖���1� H���� H��衖���UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H����: H���   H���S H���   H���S H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�W���   H�EH�UH�GH��([^_]Ð�����������SH��@A�   H��H�L$?H���  �|$? tNH�H�@�H���   H��t:H��P0���t61�H��@[�H��H��tD�Y� H�HX�K �Cu^�c�  �������H��D$,HZ�S H�ك��U �D$,��� H�HX�K �Cu�� �� H���� H�������� H����� H�����������SH��`)|$PH��o:H��H�H�HًQ ����U H�L$OA�   H���  �|$O t:H�H�P�H��B u*H���   H�L$0)|$ A�   L�D$ H��P(H�|$0�t(|$PH��H��`[Ð      �     H�H�H�HًQ ���T ��H��H��t �� H�H�H�HكI �Au7�"� ���� H�HX�K �Cu�� �� H����� H��� ����{� H����� H�����������������WVSH��PH�H��H�H�H��D��HًQ �����S H�L$OA�   H����	  �|$O t8H�H�P�H��B u(H���   H�L$0A��I��H��D$    �P H�|$0�tH��H��P[^_�H�H�H�HًQ ���S ��H��H��t �	� H�H�p�HރN �Fu7�� ���� H�HX�K �Cu�� �~� H����� H�������i� H����� H���ْ�����������VSH��XA�   H�����H��H���A    H�L$O��  �|$O tBH�H�P�H��B u2H���   H�L$0A�   E1�H��D$    �P H�D$0H��D$8�CH��H��X[^�H��H��t�� H�Hp�N �Fu7�� ����� H�Hp�N �Fu�� �� H����� H��������x� H����� H��������������SH��0H�H��H�A    H�H�HًQ �����Q H�L$/A�   H����  �|$/ t(H�H�H�H�H���   H��t9H�PH9PsH��H�PH��H��0[�L� �����H��A�PX���u�H�H�H�HًQ ���Q H��H��0[�H��H��u� � H�HX�K �Ct#�� ��� H�H�P�HڃJ �Bt�|� �w� H����� H��������� �d���H����� H���͐���������������SH��0A�   H��H�A    H�L$/H����  �|$/ t)H�H�@�H���   H�AH9A�      vH��H�AH�C   H��H��0[�@ H��PP���u�H�H�H�HًQ ���P H��H��0[�H��H��u��� H�HX�K �Ct#�� ��� H�H�P�HڃJ �Bt�u� �p� H����� H���������� �i���H���� H���Ə��������AVAUATUWVSH��0H��H��H���$  H�A    A�   H��H�L$/��  H����   �l$/@����   H�H�@�H���   H�GH9G�s  � H�SE1�I��������I�       �D  H9�~M�����   L�GH��H�GH)�M��I)�L9�IO�H����   H�H�I9�H�GH�S��   H9�� �L9��  ���tL�kA��H�       ��E��tH��������H�CH�H�H�HًQ ����N D  H��H��0[^_]A\A]A^�����H��0[^_]A\A]A^�f.�     H��������H9�t�E��t�H�C�fD  H��I9�H�Sv5H��H�GL9�s� H�S�����f.�     H�H���PHH�S�����H�H���PP���t�H�GL�G�fD  H�H���PH����E��tL�s���0�������H��H��u�}� H�HX�K �Ct#�� �b� H�H�x�H߃O �Gt��� ��� H���\� H���d����O� H�������H���?� H���G����������AWAVAUATUWVSH��XA���H��H��D����  H�A    A�   H��H�L$O�B  H���i  D�l$OE���Z  H�@�l$?H�@�L���   I�D$I9D$�)  � H�{E1�I�       �f�H9���   ����.  9���   M�\$I��M�T$I�      )�L��L)�I9�LO�I���1  �T$?M��L��L�\$0L�L$(L�T$ �`4��L�T$ L�L$(H��L�\$0L)�H��LE�M�L�M9�M�T$H�{�l  H9�A��h���H��������H9���  �����   9���   L�{E��H�       ��%���D  H��������H9��n  E����   H��H�{I�D$I;D$�0  H��I�D$ H��H��X[^_]A\A]A^A_�������D  H��������H9�tQE��tH�CH�H�H�HًQ ���K H���H��M9�H�{��   I��M�T$M9�soA�H�{�b���f�E��t�H��������H�C�E��t%fD  H��������H�{���t�9��E���H�{H��������H9���������f�     I�$L���PHH�{�����I�$L���PH�����I�$L���PP�������M�T$M�\$�H���I�$L���PP�����E���d����m���E���V����l���H��H��u�� H�HX�K �Ct#�� ��� H�H�x�H߃O �Gt�� �z� H����� H��������� H���P���H����� H���͉���������������UWVSH��(D��L�H��� H��I�H�HыQ ����   H���   H����   H���  L�I�H�H�@���  �A�  H���   H�FH9F�M  H���   � H���t  H�U0���B u2�  �     H��H�FH9���   � H�U0���B ��   H�FH�VH9�r�H�H���PP����	  H�HX�H�ًQ ����H��([^_]��H @��u
�A�K����H��([^_]�H��H����   �_��       H�H�p�HރN �F��   �b� H�HX�H���     �Q ��t���H��([^_]�H f�     H�H���PH����"����M���f�     L�IX�S H�م��^����:���fD  H�H���PHL�I�H�H�H���   H��t������������H�FH�V������k �� H�HX�K �Ct�&� �!� H���� H��葇���� H���t� H���|���������������UWVSH��(D��L�H��� H��I�H�HыQ ����   H���   H����   H���/  L�I�H�H�@���  �A�  H���   H�FH9F�M  H���   � H���t  H�U0���B u2�  �     H��H�FH9���   � H�U0���B ��   H�FH�VH9�r�H�H���PP����	  H�HX�H�ًQ ����H��([^_]�F @��u
�A�K����H��([^_]�H��H����   �� H�H�p�HރN �F��   �� H�HX�H���     �Q ��t���H��([^_]�9F f�     H�H���PH����"����M���f�     L�IX�S H�م��^����:���fD  H�H���PHL�I�H�H�H���   H��t������������H�FH�V�����i �<� H�HX�K �Ct��� ��� H���9� H���A����� H���$� H���,���������������WVSH��0H�H�@�H��H��H���   H��t_�{8 tD�KCH��H��H��0[^_�R   f�H��L�D$(�!��H�A�
   H��#��L�D$(H�@0H9�t��
   H����L�D$(D�����h ����      ��������AWAVAUATUWVSH��HH��H�A    I��M��H�L$?A�   H��E��E�������|$? ��   A�ƉD$(H�E H�@�H���   H�GH9G��  � H�uA�ωL$,H�VL9���   ����C  9D$(L�wL��  L��L��H)�L)�H��H9�HO�H���/  �T$,I��L����+��H����   H��L)���   H�I�I9�H�GH�u�2  H�V� L9��y��������  9D$(��  M���Z  A�$ �   � H�H���PP�M��~kA�$ H�} uh�   H�E H�H�H�Q �gC �NL��H��H����  �� H�E H�p�H�N �F��  �� M����  f�     H�UH��t�H��H��H[^_]A\A]A^A_� I��L��L���*��H�GH�uL�wH������A�$H�GI�\$H�WH�EH9�sCH��H�GH9�sv� I��H�u�Q����    H�H���PHH�u�8���H�H���PH����H�H���PP�����   M��~� H�u�   H���������������   ��D  H�H���PHH�uI�������L�wL� M9�H�U�y���M�OM��L�O�w��������L���M��~�A�$ H�}҃����b���H�GH�W�����h����U� H�E Hh�M �Et7��� ��� � H�} ��������H���>� H���F������������� H���� H���'����������VSH��8H�H��H�A    H�H��HًQ ����8A H�L$/A�   H���%����|$/ t.H�H�H�H�H���   H��tEH�HH9Hs@:q�uH��H�HH��H��8[^�fD  �      L� @��H��A�PX���u�H�H�H�HًQ ���@ H��H��8[^�H��H��u�0� H�HX�K �Ct#��� �� H�H�p�HރN �Ft�� �� H���� H�������� �]���H����� H�������������������WVSH��0H��H�A    H��L��H�L$/A�   H�������|$/ ttH�H�@�H���   H�AH+AtgH��~mH�H9�HN�I��H�R�H���   H��L�	A�Q@H�CH��0[^_�H��H��tR�3� H�H�x�H߃O �Gui�:� H�CH��0[^_�H��P8H���H���u�H�H�H�HًQ ���X? ���� H�HX�K �Ct�{� �v� H���޻ H����~���a� H���ɻ H����~���UWVSH��(H�iH��H��H���- 1�H��Hǃ�       f���   H��� H�H��(H�CH�GHǃ�       Hǃ       Hǃ      H�CH�Hǃ      H�p�H�H���g! H���   H���h; H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H�G    H��([^_]�H��H�OK H��H�PH�S�O- H����}���������WVSH�� H�qH��H��H���w, 1�H��H��f���   H�y� H�H��(Hǃ�       Hǃ�       Hǃ       Hǃ      Hǃ      H�CH�C    �; �H�� [^_�H��H��J H��H�PH�S�, H���}���������WVSH�� H�qH��H����+ 1�1�H��f���   H�͸ H�H��(Hǃ�       Hǃ�       Hǃ       Hǃ      Hǃ     �       H�CH�C    �; �H�� [^_�H��H��I H��H�PH�S��+ H���k|�������������WVSH�� H�L��H�L�BH�P�L�H�WH�QHH�H�H��H�p�H�H���C H���   H���D9 H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H�G    H�� [^_Ð�����H�H�L�JH�P�L�L��H�A    HH��
: ����������H�H�L�BH�P�L�1�H�A    HH���9 �����������SH�� H�<� H�H��H H��H�A    H�IH��H��* H��H�� [鲳 ��H�� H�H�H H��H�A�    H��H��w* �������H�H�H�@�H�RH�H�A    Ð����UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���� H���   H����7 H���   H���7 H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�U���   H�GH�WH�EH��H��([^_]Ð��������H�␐�����������SH�� H�H��H�H�H���H��H�� [Ð��SH�� H�H��H�H�H���H��H�� [Ð��VSH��8E1�H��H��H�L$.H��������|$. tBH�H�H�H�H��tBH���   L�D$/H����c H���T$/t@��tH��   H�H�H��H��t=H��H��8[^ú   Q �9 H��H��8[^�D  H�H�H�Hـ�҃������H��   H�H�H���H��H��t �ʳ H�H�p�HރN �Fu7�ѵ �誳 H�HX�K �Cu�D� �?� H��觵 H���x��      ��*� H��蒵 H���x�������������K�������������������������������������������������������������K��������������VSH��   E1�H��H��H�L$wH���a����|$w ��   H��D$x    H�P�H�H��H��   H����   L�H�L$`A�����L���   L�D$XL�D$HL�D$|L�D$0L�D$xL�D$(L�D$PL�L$PL�L$@H�D$@    H�D$ A�R�D$|��T$x��uH��H�Ĉ   [^�f�H�H�H�H�Q �7 H��H�Ĉ   [^��[ H��H��t �� H�H�p�HރN �Fu7�%� ���� H�HX�K �Cu蘸 蓸 H����� H���w���~� H���� H����v�����������������+���������������k�����������������������������VSH��   E1�H��H��H�L$wH��������|$w ��   H��D$x    H�H�H�H��   H��H����   L���   A�����H�D$@    L�L�D$XH�L$`L�D$HL�D$|L�D$0L�D$xL�L$PL�L$@L�D$(L�D$PH�D$ A�R�D$|�T$x= ���} ��� ����T$xf���u'H��H�Ĉ   [^�=�  ~7����  �҉T$xf�t�H�H�H�H�Q ��5 H��H�Ĉ   [^�D  f����Y H��H��t'�X� H�H�p�HރN �Fu>�_� �T$x�w����1� H�HX�K �Cu�˶ �ƶ H���.� H���6u��豶 H���� H���!u����[���������������������������������������������WVSH��0H�\$ H�Ή�H��H���  �|$  t!H�H�@�H���   H�A(H;�      A0sH@�8H�A(H�D$(H�HB��@ H��t �Z ��uH���   H��tH��P0���t7H��H��0[^_�H�@���Ph���u�H�H�H�H�Q ���4 �fD  H�L$(H�HH�Q ���i4 �H��H���  H���t��H��H��u�֮ H�Hp�N �Ft-�p� 軮 H�H�x�H��O �Gt�R� 轰 �����C� H��諰 �H��衰 닐��������������VSH��(H�HH�H�H��H�X�H�H���� H���   H���0 H���   H���0 H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   ���   H��([^Ð��������SH�� H�H�@�H��H���   H��tH��P0���t	H��H�� [�H�H�H�HًQ ����2 H��H�� [�H��H��t �t� H�H�P�HڃJ �Bu7�{� ��T� H�HX�K �Cu�� �� H���Q� H���Yr���Գ H���<� H���Dr������SH��@H�L�
L�RH��H�H�H��A u/H���   L�D$ L�L$ A�   H�L$0L�T$(H��P(H�|$0�tH��H��@[�f�     H�H�H�HًQ ���2 H��H��@[�H��H��t 脬 H�H�P�HڃJ �Bu7苮 ��d� H�HX�K �Cu��� ��� H���a� H���iq���� H���L� H���Tq������SH��@H�H��H�H�H��A u,H���   H�L$0E��I��L�H���D$    A�R H�|$0�tH��H��@[� H�H�H�HًQ ���+1 H��H��@[�H��H��t 褫 H�H�P�HڃJ �Bu7�      諭 �脫 H�HX�K �Cu�� �� H��聭 H���p���� H���l� H���tp������VSH��HH�H��H�����H���A    H�H�H��A u2H���   A�   E1�H�L$0H��D$    �P H�D$0H��D$8�CH��H��H[^�H��H��t�̪ H�Hp�N �Fu7�֬ ��诪 H�Hp�N �Fu�I� �D� H��謬 H���o���/� H��藬 H���o�����������������UWVSH��8H�\$ H��H��H��H��L���/  �|$  t H�I��H��H�@�H���   H��P`H9�uHH�D$(H�HB��@ H��t �T ��uH���   H��tH��P0���t3H��H��8[^_]��    H�H�H�H�Q ���+/ �f�     H�L$(H�HH�Q ���	/ �H��H��u艩 H�Hp�N �Ft#�#� �n� H�H�x�H��O �Gt"�� � � H���h� H���  H���hn���S� ����H����H���A� �א��������������SH��0H�H��� H�QH�H�H�H��H���   D�@ H��t5E��tD��H����H��0[�<. H�T$(�����H�T$(H�HP�D�B H��E��u��H��0[ÐSH��0H�H��� H�QH�H�H�H��H���   D�@ H��t5E��tD��H����H��0[��- H�T$(����H�T$(H�HP�D�B H��E��u��H��0[ÐVSH��(H�AH�H��HB��@ H��t �R ��uH���   H��tH��P0���tH��([^�H�NH�HH�Q ��H��([^�@- VSH��(H�AH�H��HB��@ H��t �^R ��uH���   H��tH��P0�      ���tH��([^�H�NH�HH�Q ��H��([^��, VSH��(H�H�@�H��L��H���   H��P`H9�u
H��([^� H�HX�S H�ك�H��([^�, �����AUATUWVSH��hH�l$PH��I��H��H��������|$P ��   H�H�X�H�H���   H���U  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D�D$ L�D$0L�d$(�PH�|$H tH�H�H�H�Q ����+ H�D$XH�HB��@ H��t$�Q ��uH���   H��tH��P0�����   H��H��h[^_]A\A]� L���   M����   A�}8 t)E�EYD�����   H�ƃ�   H�X�H��!���D  L�����I�E H��	��A�    L�H0�    I9�t��    L��A��D����     H�L$XH�HH�Q ����* �Q�����N ��N H��H��u.�l� H�Hp�N �Ft6�� H��H������H���sj���>� H�H�x�H��O �Gt�ի �Ы H���8� ���1� ����H���$� 믐�AUATUWVSH��hL�d$PH�Ή�H��L��������|$P ��   H�H�X�H�H���   H���G  ���    @����   ���   L���   H�L$@�    I��M��L�D$0L�D$0��H�D$8H�E �T$ H��|$(�P�|$H tH�H�H�H�Q ���) H�D$XH�HB��@ H��t$��N ��uH���   H��tH��P0�����   H��H��h[^_]A\A]�f�L���   M����   A�}8 t)A�UY�Ј��   H�ƃ�   H�X�H��$���fD  L�����I�E H�����    L�@0�   �       I9�t�L��A�����H�L$XH�HH�Q ����( �a�����L ��L H��H��u.�[� H�Hp�N �Ft6��� H��L���
���H���bh���-� H�H�x�H��O �Gt�ĩ 迩 H���'� ��� � ����H���� 믐ATUWVSH��p)t$`H�l$PH��H��H��f(������|$P ��   H�H�X�H�H���   H���Q  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D�D$ L�D$0�t$(�P8�|$H tH�H�H�H�Q ���' H�D$XH�HB��@ H��t$��L ��uH���   H��tH��P0�����   (t$`H��H��p[^_]A\�L���   M����   A�|$8 t%E�D$YD�����   H�ƃ�   H�X�H�����L�����I�$H����A�    L�H0�    I9�t��    L��A��D���fD  H�L$XH�HH�Q ����& �V����J �J H��H��u.�<� H�Hp�N �Ft6�֧ H��H�������H���Cf���� H�H�x�H��O �Gt襧 蠧 H���� ���� ����H����� 믐�ATUWVSH�Ā�*�|$0H�l$pH��H��H�������|$p ��   H�H�X�H�H���   H���d  ���    ��   D���   H���   �    I���l$0H�L$`H��H�T$P�|$@H�T$@��H�D$XH�H�T$(H��D�D$ L�D$P�P@�|$h tH�H�H�H�Q ���~% H�D$xH�HB��@ H��t$�J ��uH���   H��tH��P0�����   H��H��[^_]A\��    L���   M����   A�|$8 t(�      E�D$YD�����   H�ƃ�   H�X�H����� L���X��I�$H����A�    L�H0�    I9�t��    L��A��D����     H�L$xH�HH�Q ���$ �O����H �zH H��H��u.�� H�Hp�N �Ft6覥 H��H������H���d���ޞ H�H�x�H��O �Gt�u� �p� H���ؠ ���Ѡ ����H���Ġ 믐�AUATUWVSH��hH�l$PH��A��H��H���n����|$P ��   H�H�X�H�H���   H���U  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D�D$ L�D$0D�d$(�P�|$H tH�H�H�H�Q ���\# H�D$XH�HB��@ H��t$�H ��uH���   H��tH��P0�����   H��H��h[^_]A\A]� L���   M����   A�}8 t)E�EYD�����   H�ƃ�   H�X�H��!���D  L���8���I�E H�m��A�    L�H0�    I9�t��    L��A��D����     H�L$XH�HH�Q ���y" �Q����_F �ZF H��H��u.�� H�Hp�N �Ft6膣 H��H������H����a��辜 H�H�x�H��O �Gt�U� �P� H��踞 ��豞 ����H��褞 믐�AUATUWVSH��hH�l$PH��A��H��H���N����|$P ��   H�H�X�H�H���   H���U  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D�D$ L�D$0D�d$(�P �|$H tH�H�H�H�Q ���<! H�D$XH�HB��@ H��t$�bF ���      uH���   H��tH��P0�����   H��H��h[^_]A\A]� L���   M����   A�}8 t)E�EYD�����   H�ƃ�   H�X�H��!���D  L������I�E H�M���A�    L�H0�    I9�t��    L��A��D����     H�L$XH�HH�Q ���Y  �Q����?D �:D H��H��u.�̚ H�Hp�N �Ft6�f� H��H���{���H����_��螚 H�H�x�H��O �Gt�5� �0� H��蘜 ��葜 ����H��脜 믐�AUATUWVSH��hH�l$PH��I��H��H���.����|$P ��   H�H�X�H�H���   H���U  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D�D$ L�D$0L�d$(�P(�|$H tH�H�H�H�Q ��� H�D$XH�HB��@ H��t$�BD ��uH���   H��tH��P0�����   H��H��h[^_]A\A]� L���   M����   A�}8 t)E�EYD�����   H�ƃ�   H�X�H��!���D  L�������I�E H�-���A�    L�H0�    I9�t��    L��A��D����     H�L$XH�HH�Q ���9 �Q����B �B H��H��u.謘 H�Hp�N �Ft6�F� H��H���[���H���]���~� H�H�x�H��O �Gt�� �� H���x� ���q� ����H���d� 믐�AUATUWVSH��hH�l$PH��I��H��H�������|$P ��   H�H�X�H�H���   H���U  ���    ��   D���   H���   H�L$@�    I��H��H�T$0H����H�D$8H�D��      D$ L�D$0L�d$(�P0�|$H tH�H�H�H�Q ���� H�D$XH�HB��@ H��t$�"B ��uH���   H��tH��P0�����   H��H��h[^_]A\A]� L���   M����   A�}8 t)E�EYD�����   H�ƃ�   H�X�H��!���D  L�������I�E H����A�    L�H0�    I9�t��    L��A��D����     H�L$XH�HH�Q ��� �Q�����? ��? H��H��u.茖 H�Hp�N �Ft6�&� H��H���;���H���[���^� H�H�x�H��O �Gt��� �� H���X� ���Q� ����H���D� 믐�WVSH�� H�yH��H��H���
 1�H��Hǃ�       f���   H�Q� H�H��(H�CH�Hǃ�       Hǃ�       Hǃ       Hǃ      Hp�H����� H���   H���� H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H�� [^_�H��H��' H��H�PH�S��	 H���\Z��������������WVSH�� H�qH��H��H���	 1�H��H��f���   H�Y� H�H��(Hǃ�       Hǃ�       Hǃ�       Hǃ       Hǃ      H�C�J �H�� [^_�H��H�7' H��H�PH�S�7	 H���Y�����������������SH�� H��H�I�_ 1�Hǃ�       f���   H��� H�H��(Hǃ�       Hǃ�       Hǃ       Hǃ      H�CH�� [Ð������WVSH�� H�qH��H���� 1�1�H��f���   H�=� H�H��(Hǃ�       Hǃ�      �       Hǃ�       Hǃ       Hǃ      H�C�. �H�� [^_�H��H�& H��H�PH�S� H���X�����VSH��(H�H�HH�H�BH��H�I� H�p�L�H���� H���   H��� H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H��([^�L�
L�	II�H�BL��H��g �������H�H�H�@�H�RH�Ð������������H�H�HH�H�B1�H��( ��������SH�� H�ܓ H�H�
% H��H�IH��H�� H��H�� [�
� ����������H��� H�H��$ H��H��H��� ���������������H�H�H�@�H�RH�Ð������������WVSH�� H�H�p�H��H�H�H�X�H��H�H���G� H���   H��� H���   H���	 H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   ���   H��H�� [^_Ð�������������H�␐�����������SH�� H�H��H�H�H���H��H�� [Ð��SH�� H�H��H�H�H���H��H�� [Ð������������������WVSH��@H�|$0H��H��H��H�������|$0 t<H�H�H�H�H��trH���   L�D$/H���9@ H��uH��   H�H�H��M H��thH�D$8H�HB��@ H��t �; ��uH���   H��tH��P0���tH��H��@[^_ú   Q � �H�L$8H�HH�Q ��� ��H��   H�H�H���H��H�������H���U��H��H��u�� H�Hp�N �Ft-�{� �Ə�       H�H�X�H�K �Ct�]� �ȑ �(����N� H��趑 �H��謑 닐������������x������������{��������������H��8�*�|$ H�T$ �|���H��8Ð�������Z��G�����������������������������������������k���������������{��������������H�H�@�D��J��@t��t���0������(��������������8������������K���������������[������������������H)�H������@H��   �M�ÐH�Ð�����������H�Ð�����������SH�� H��@�H�˅�~E1�E1�1���  H��@�����H�� [ÐWVSH�� H�ˉ�1��-  H��L�HH��tH��t,L��@��I������I��L���F    H��D H�� [^_�@�x�����������WVSH�� H)�H��H��1�H����  H��L�HH��t<H��u$L���F    H��D H�� [^_�f.�     L��I��H������I������F�������WVSH�� H��H��tH��tWH)�H��1�H���L  H��L�HH��t2H��uL���F    H��D H�� [^_�L��I��H���"���I������F��H�� �: ���������WVSH�� H��H��tH��tWH)�H��1�H����  H��L�HH��t2H��uL���F    H��D H�� [^_�L��I��H������I������F��H��� �9 ���������H�)� Ð�������I)�I��tM��uÐ�[�����Ð����I)�I��tM��uÐ�;�����Ð����I)�I��tM��uÐ������Ð����I)�I��tM��uÐ�      �������Ð����H��(H�H�P�H9P�rH��(�f.�     1��Y  �H��(�H��苋 �H��(額 �UWVSH��(H��������?�l$pH��H�L�H��L��H+B�I9�wAH����  H��tH>H��H��t@��I���M���H��H��([^_]ÐH��@�/H��([^_]�H��� �U9 �����UWVSH��(H�\$pL��I��H��H���  H��tH>H��H��t!I��H�������H��H��([^_]�f.�     �E �H��H��([^_]Ð����������������h�����������VSH��(H�L�@�H��H��L9�s�P���x����H�H�H��([^�H�P� ��> ���SH�� H��P�H�˅�x�����H�H@�H�� [Ð������������ˇ ������������������A��~Ð髇 �������������AH�AÐ�����H�AÐ����������H��� Ð��������A����Ð��������A    Ð��������A    H��D �D�AH�AE��x�� H�A�f.�     E1��   ��������VSH��(H��H�	L�I��H�V�U   L�L�HH��M��tI��t0H�VL���D���L�I��L���C    L�B�D H��([^�@ �F�CL��֐���SH�� H��������?H9�H��wWH�IH9�v8H�H9�HB�H�K9H��   vH9�sH��   ���  H)�H9�HG�H�K胆 H�X�@    H�� [�H��� �6 ������VSH��(H�H��H�H�P�H�Y���xH�������H�H�H��([^�VSH��(H��H�
H�֋A���xH�������H�H��H�H��([^Ð�H�D�@�E��y�@�    L�E�H�E��yA�@�    L�      �H�Ð�SH�� H��P�H�˅�x�i���H�H�� [�E1�1�H�L�@��O  ���������������VSH��(E1�A�   H��H+H��H���   H��@�����H�H��([^Ð�����������VSH��(I)�H��H��uH��([^��     H+E1�H��H����  H��@�����H�H��([^Ð����������SH�� H�L�H�H��L��H)�L9�LF�L9�wE1�H���  H��H�� [�H��� I��H�G� �5; �����SH�� H��P�H�˅�x�I���H�H�� [�VSH��(H��H��H���<���H��H��I��H��([^�   ��������WVSH�� M��H��H��twH��������?H�H�p�H)�I9���   L�H;p���   H9�wH�P�H�H9�vGH��H��L�D$P��  H�L�D$PHI�I��tMH������H��@�    H�p��0 H��H�� [^_�H��H��H)�L�D$P�y  H�L�D$PH�HI�I��u���봋@���~H��j���H�	�H��� ��3 �������������UWVSH��(H�H�p�H��H��H��tEH�H�h�H�H;h�vFH��H����  H�H�HI�H��tBI���S���H��@�    H�h��( H��H��([^_]�D  �@����H�H�HI�H��u���뿐�UWVSH��(H�H�X�H��H��I9�w}L)�L9�IG�H��tYH�H�h�H�H9h�r�@���~H��H��L�D$`�P  L�D$`H�H�L�HI�H��t(I������H��@�    H�h��( H��H��([^_]�f�����H�@� I��H�� �8 ���H��H�L�@������SH�� H��H��t	E���
   H��H�� [ÐUWVSH��(H��������?H��H�	H��D��H��      Y�H)�H9�raH�H;Y�v?H��H���
  H�HI�H��t;@��I�������H��@�    H�X�� H��([^_]ËA����H�HI�H��u�@�)��H�l� �1 ���������H��(�W���H��H��(Ð��������������VSH��(H��H��H�������H��H��I��H��([^�   ��������VSH��8H�L��I��H��L�@�H��������?H9���   L9�vH�t$ 1�H�������H��8[^�J� I9�w�@���~H�L�@��� H�	L��H)�H9�v6H��tH��tGI��L������H�f�     �A�    H��H�q��1 �H��tH��t�I��L������H��ѐA��H���H�'� �0 ���������VSH��8H�2H91H��t'�V�H�N�H�A��x"�� H��������A���~H�3H��H��8[^�H�T$/E1�����H����H��� �֐H��(H�L�R�L��L)�L9�IG�M9�wL�I��H��(����H��� M��H�c� �6 ��������������H��H�L�@�a����H��8H�H�@�E��I��1�D�D$ I�������H��8Ð���������M�HH+M� �   �VSH��8A�   H��H+E��H��D�D$ E1�H������H��@�����H�H��8[^Ð��H��8H+E��D�L$ M��E1��U����H��8Ð��������������WVSH�� H��L��H��L���h���I��H��H��I��H�� [^_�    UWVSH��8H��H�L��H��L�J�L9��5  H��������?L)�H9��  L9�v$M��H�|$ E1�H��H���>���H��8[^_]�D  I�M9�wԋB����L��I��E1�H+1H���  L�I�1I�H�:L9�wH��t}H��tpI��L���      ���H���L9�r!H��tsH��tPI��H��L�������H���{���H)�H��tGH��tL��I�������I��I�9I��I�)I)�I��t6M��t����H���9����A�H���+����A���� A�H��������H������H��� �- H��� I��H��� �3 ����M� M�H���������H��(M�L�T$PM�C�L��M��I)�M9�MG�L9�wM�H��(�N���H��� M��I��H��� �E3 �����H��8H�H�@�E��H9�wD�L$ M��E1�����H��8�H�`� I��I��H�A� ��2 ��������������VSH��(H��H�
H�֋A���xH������H�HI�H��H�H��([^Ð�������������E1��   ��������H��(I��������?H�L9�H�@�w8H9�w#rH��(�f.�     H)�E1�I��H��(�  H)�E��H��(�����H��� �, ��I��tM��u�@ �������Ð����H��H�Ð��������H��@���y�D  �+��������������I��tM��u�@ ������Ð����L)L$(H��H+I)��  �������������UWVSH��8H��H��L��L��L�������H��H+I��H�D$ I��I)�H���H  H��8[^_]Ð��������������L)L$(H��H+I)��  �������������H��H+I)��  ��H��8M�	M�Q�H��H+I)�L�T$ ��   H��8Ð������������L)L$(H��H+I)��   �������������L)L$(H��H+I)��   �������������H��8M�QH��L�T$ H+M�	I)��r   H��8Ð������������D�T$(H��H+D�T$(I)��w�����������      UWVSH��8H��L��H��L��L������I��I��H��H�D$ H���   H��8[^_]Ð����AUATUWVSH��HH��$�   H��L��H��H�L�H�L9��-  L��H)�H��������?L9�IG�L)�H�H9��  H9�v)I��H�l$ H��I��H���B���H��H��H��H[^_]A\A]�I�I9�rϋ@����H�H�)L�8L9���   L�I�L9�r@H)�H�H)�I��H��H��I��I���  H�J�!H�H��tsH��t�I��������@ L�l$?E1�M���`���H�l$ I��H��I��H��I������H�Ƹ�����A�D$����A���I�L$��6x �2����H)�I���q���D  ������H�� I��H�� ��. H�� �( I�L$�H��L���$���H���L?��������������H��8M�	I�A�H�D$ �K���H��8Ð�����SH�� I�L�T$PL�\$XL�K�L��L)�L9�IG�M9�wN�H�D$PH�� [����H��� M��H�t� �. ���������������H��(H�D�\$PL�P�L��H)�L9�LF�L9�wD�\$PH��(�����H�(� I��M��H�� ��- ������SH��@H��H�	H;Q�tTH�A�H9�HB�H��I��H�T$?I)������H��������Q���~H�H��@[�fD  H��H�D$(�v H�D$(�܋A���~�H�렐��������������H��(E1�H�H�@�H�P�H9�wA�   H��(�J   H� � I���H�X� �- ���H��tH��u�@ A��I�Љ�����f�D�Ð�����������AWAVAUATUWVSH��8H�H�p�M�4I��L��H�P�L)�H��M��H�L)�H9�w�@�����   H�H�P�L�D$/H�������      M��H�xI��tH�U H�xI����   M��H�������H��H�U u6�������B���~xH�} �G�    H�_�� H��8[^_]A\A]A^A_�@ K�L,L�L�H��toI������H�U 뫐H��H�9t�M9�t�J�7M�H��J�'tRI���r���H�} �@ H�J���t �z���f��H��A�GH�U �V����f.�     ��H�U �<���f���H�} �>�����UWVSH��(H�H�x�H�ˉ�H�wH;p�w�@���~H��H������H�H�P�@�,H��@�    H�p��D8 H��([^_]Ð��������SH��0H�L�D$/H��H�1�1��T���H�H��0[Ð����������VSH��(H��H��H������H��tH��L�D$P�����L�D$PH�E1�H�������H�H��([^Ð������������SH�� L��H��E1�H��J�I������H�H�� [Ð���������SH�� H��I��1�1�����H�H�� [Ð��SH��0H�D�@�H��H�H�H�QE��x��H�H��0[��    H�T$/E1��3���H�H��0[Ð���������SH�� H��H�
L��L�I�J�	M9�wL�E1�I���w���H�H�� [�H��� H� � �) �����������SH��0H��H�
H�A�H��L)�L9�IG�L�H�I9�wL�E1�L�D$/����H�H��0[�H�+� I��H��� �J) ����������SH�� H��H�
H�A�H��L)�L9�IG�L�H�I9�wL�L�D$PE1�����H�H�� [�H�˷ I��H�?� ��( ����������SH�� E1�H�BH��H�
H�H�������H�H�� [Ð���������SH��01�L�D$/H��1������H�H��0[ÐSH�� H��H��A��M�      �������H�H�� [�SH�� H��H��L��M��E1�����H�H�� [Ð�������������SH�� H��H��L��M��E1��W���H�H�� [Ð�������������SH�� H��H��L��M��E1�����H�H�� [Ð�������������SH��0H�L�D$/H��H�1�1��$���H�H��0[Ð����������VSH��(H��H��H������H��tH��L�D$P�����L�D$PH�E1�H������H�H��([^Ð������������SH�� L��H��E1�H��J�I���s���H�H�� [Ð���������SH�� H��I��1�1��|���H�H�� [Ð��SH��0H�D�@�H��H�H�H�QE��x��H�H��0[��    H�T$/E1�����H�H��0[Ð���������SH�� H��H�
L��L�I�J�	M9�wL�E1�I���G���H�H�� [�H�Y� H�г �{& �����������SH��0H��H�
H�A�H��L)�L9�IG�L�H�I9�wL�E1�L�D$/�����H�H��0[�H��� I��H�o� �& ����������SH�� H��H�
H�A�H��L)�L9�IG�L�H�I9�wL�L�D$PE1�����H�H�� [�H��� I��H�� �% ����������SH�� E1�H�BH��H�
H�H�������H�H�� [Ð���������SH��01�L�D$/H��1������H�H��0[ÐSH�� H��H��A��M������H�H�� [�SH�� H��H��L��M��E1������H�H�� [Ð�������������SH�� H��H��L��M��E1��'���H�H�� [Ð�������������SH�� H��H��L��M��E1��w���H�H�� [Ð������������������H�	��A���~�H����m ����������H�	�      ��A���~�H���m �����H��(�����H��H��(Ð��������������VSH��(H��H��H���|���H��H��I��H��([^�������������k��������������SH�� H��H�H��L�@�i���H��H�� [�SH��0A�   H�L�@���H�ˉT$ 1������H��H��0[Ð���VSH��(H�H�֋P�H�˅�x�����H�H�H��([^Ð�������VSH��(H��H��H������H��H��I��H��([^�������������k��������������H��H�L�@�a����UWVSH��(H�H�x�H�ˉ�H�wH;p�w�@���~H��H���P���H�H�P�@�,H��@�    H�p��D8 H��H��([^_]Ð������A�%H�J��tH�J�B+��t�#H��A��A��  A��  tJH�QA�.*  E��fD�u?L�BA��tF���� @  A��   t=A��  tF����� ��G�A�  ÐE��H��t.D�H��A��L�Bu��fA�  Ã���� ��E�A�  �H��L�A% @  ����� ��A�A�  Ð��������������SH�� H�$o H��H��� �   H��H�� [�'k �������H��n H�� �H�Y� � Ð�����SH�� H�AH��H����   �@!.H�C�@",H�SH�d� H�BH�SH�B    H�SH�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H��� H�S� �B\H�S�B`H��� L� 1�f.�     A� H�S�LdH��H��u�H�� [� �p   �Vj H�O~ 1��@    H�H�@    H�@    f�P �@" H�@(    H�@0    H�@8    H�@�      @    H�@H    H�@P    H�@X    �@`    �@o H�C��������������������VSH��(1�M��H�QH����E1�1҉AH��m H��t����H��([^�H��H���a# H���0�����������VSH��(1�M��H�A    H�����AH�=m H��%����H��([^�H��H���# H���j0������������VSH��(1�H��H�A    H����E1�1҉AH��l H�������H��([^�H��H���" H���0�������VSH��(1�M��H�QH����E1�1҉AH��l H������H��([^�H��H���q" H����/�����������VSH��(1�M��H�A    H�����AH�Ml H��5����H��([^�H��H���"" H���z/������������VSH��(1�H��H�A    H����E1�1҉AH��k H�������H��([^�H��H����! H���%/�������VSH��(H���"   H��H��([^�g H��H���g H����.���VSH��(H�� H��H��H�H�IH��tH��PH��H��([^�\! H��H���Q! H���.�����������SH�� H�AH��H����   �@!.H�C�@",H�SH��� H�BH�SH�B    H�SH�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�� H�S� �B\H�S�B`H��� L� 1�f.�     A� H�S�LdH��H��u�H�� [� �p   �f H��z 1��@    H�H�@    H�@    f�P �@" H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@o H�C�������������      ��������VSH��(1�M��H�QH����E1�1҉AH�<j H��t����H��([^�H��H��� H����,�����������VSH��(1�M��H�A    H�����AH��i H��%����H��([^�H��H���R H���,������������VSH��(1�H��H�A    H����E1�1҉AH��i H�������H��([^�H��H���� H���U,�������VSH��(1�M��H�QH����E1�1҉AH�Li H������H��([^�H��H��� H���	,�����������VSH��(1�M��H�A    H�����AH��h H��5����H��([^�H��H���b H���+������������VSH��(1�H��H�A    H����E1�1҉AH��h H�������H��([^�H��H��� H���e+�������VSH��(H���"   H��H��([^��c H��H����c H���1+���VSH��(H�S� H��H��H�H�IH��tH��PH��H��([^� H��H��� H����*�����������SH�� H�AH��H����   �.   �,   f�P"H�Cf�H$H�CH�ڥ H�HH�CH�@    H�SH��� H�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�5� H�S� �B\H�S�B`H�.� L� 1�f�     fA� H�Sf�LBdH��H��u�H�� [Ð��   ��b H��v �@    H�H�@    H�@    �@  �@"    H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@z H�C������������������VSH��(1�M��H�QH����E1�1҉AH��      �f H��d����H��([^�H��H���� H���))�����������VSH��(1�M��H�A    H�����AH��f H������H��([^�H��H��� H����(������������VSH��(1�H��H�A    H����E1�1҉AH�8f H�������H��([^�H��H���- H���(�������VSH��(1�M��H�QH����E1�1҉AH��e H��t����H��([^�H��H���� H���9(�����������VSH��(1�M��H�A    H�����AH��e H��%����H��([^�H��H��� H����'������������VSH��(1�H��H�A    H����E1�1҉AH�He H�������H��([^�H��H���= H���'�������VSH��(H���"   H��H��([^�` H��H����_ H���a'���VSH��(H��� H��H��H�H�IH��tH��PH��H��([^�� H��H���� H���'�����������SH�� H�AH��H����   �.   �,   f�P"H�Cf�H$H�CH�
� H�HH�CH�@    H�SH�� H�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�e� H�S� �B\H�S�B`H�^� L� 1�f�     fA� H�Sf�LBdH��H��u�H�� [Ð��   ��^ H�Os �@    H�H�@    H�@    �@  �@"    H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@z H�C������������������VSH��(1�M��H�QH����E1�1҉AH�|c H��d����H��([^�H��H��� H���Y%����      ��������VSH��(1�M��H�A    H�����AH�-c H������H��([^�H��H��� H���
%������������VSH��(1�H��H�A    H����E1�1҉AH��b H�������H��([^�H��H���] H���$�������VSH��(1�M��H�QH����E1�1҉AH��b H��t����H��([^�H��H��� H���i$�����������VSH��(1�M��H�A    H�����AH�=b H��%����H��([^�H��H���� H���$������������VSH��(1�H��H�A    H����E1�1҉AH��a H�������H��([^�H��H���m H����#�������VSH��(H���"   H��H��([^�4\ H��H���)\ H���#���VSH��(H��� H��H��H�H�IH��tH��PH��H��([^�� H��H���� H���I#�����������SH�� H�AH��H���K  H�7� H�3� H�H@H�XHH�'� H�'� H�HXH�X`H�� H� � H�HhH�XpH�� H�� H�HxH�ж H���   H�� H�PH�	� H�PH���   H��� H���   H�� H�� H�P H�P(H��� H���   H�Ѷ H���   H�˶ H�P0H�P8H�PPH��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H�{� H���   H�_� H���   H�f� H��   H�b� H���   H��  H�U� H��  H�P� H��H  H�[� H��P  H�Q� H��X  H�G� H��  H�!�      � H��`  H�/� H��   H�	� H��(  H��� H��h  H�	� H��0  H�� H��8  H�� H��p  H�� H��@  H��x  H���  H�� [ù�  �Y H��� �@    H�@    H�@    H�QH�@     H�H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    H�@`    H�@h    H�@p    H�@x    Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ       Hǀ      Hǀ      Hǀ      Hǀ       Hǀ(      Hǀ0      Hǀ8      Hǀ@      HǀH      HǀP      HǀX      Hǀ`      Hǀh      Hǀp      Hǀx      Hǀ�      ƀ�   H�C����������VSH��(1�M��H�QH�����AH�!] H��i 1�H��H�C �[����H��([^�H��H���( H���������������������ATUWVSH�� 1�M��H�A    L��H����H�ՉAH��\ H��� H��H��H���������uH�s H��H��������H�� [^_]A\�H������L�`L���V M��H��H�������H�C ��H��H���{ H������H���X H�K H9�t
H��t�8V �3_ H���Z �Ɛ��������VSH��(1�H��H�A    H�����AH��[ H��5 1�H��H�C �'���      ��H��([^�H��H���� H���L��������������VSH��(1�M��H�QH�����AH��[ H��� 1�H��H�C ������H��([^�H��H��� H����������������������ATUWVSH�� 1�M��H�A    L��H����H�ՉAH�#[ H��k H��H��H���M�����uH�s H��H���J����H�� [^_]A\�H������L�`L���U M��H��H���\���H�C ��H��H���� H���C��H���W H�K H9�t
H��t�T �] H���Y �Ɛ��������VSH��(1�H��H�A    H�����AH�]Z H�� 1�H��H�C �����H��([^�H��H���d H�����������������SH�� H���   H��H�� [�&T ������VSH��(H��Y H�q H�H���4 H9�tH��tH����S H�KH��tH��PH�K� H��H��([^�� ������������VSH��(H��Y H�q H�H���� H9�tH��tH���S H�KH��tH��PH�K�Z H��H��([^�| ������������SH�� H�AH��H���K  H�ʯ H�ɯ H�H@H�XHH��� H�ǯ H�HXH�X`H�Ư H�ϯ H�HhH�XpH�ԯ H�߯ H�HxH�P� H���   H�ԯ H�PH�ۯ H�PH���   H�7� H���   H�ï H�į H�P H�P(H�%� H���   H��� H���   H��� H�P0H�P8H�PPH��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H���   H��� H��      ��   H�j� H���   H��� H��   H��� H���   H��  H��� H��  H��� H��H  H��� H��P  H��� H��X  H��� H��  H�e� H��`  H��� H��   H�Q� H��(  H�K� H��h  H�m� H��0  H�7� H��8  H�Y� H��p  H�S� H��@  H��x  H���  H�� [ù�  �6Q H�/� �@    H�@    H�@    H�QH�@     H�H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    H�@`    H�@h    H�@p    H�@x    Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ�       Hǀ       Hǀ      Hǀ      Hǀ      Hǀ       Hǀ(      Hǀ0      Hǀ8      Hǀ@      HǀH      HǀP      HǀX      Hǀ`      Hǀh      Hǀp      Hǀx      Hǀ�      ƀ�   H�C����������VSH��(1�M��H�QH�����AH��T H��� 1�H��H�C �[����H��([^�H��H��� H���������������������ATUWVSH�� 1�M��H�A    L��H����H�ՉAH�cT H�� H��H��H���m�����uH�s H��H��������H�� [^_]A\�H���&���L�`L���:N M��H��H���|���H�C �      ��H��H��� H���c��H���+P H�K H9�t
H��t��M ��V H���+R �Ɛ��������VSH��(1�H��H�A    H�����AH��S H��� 1�H��H�C �'����H��([^�H��H��� H������������������VSH��(1�M��H�QH�����AH�AS H��i 1�H��H�C ������H��([^�H��H���( H���������������������ATUWVSH�� 1�M��H�A    L��H����H�ՉAH��R H��� H��H��H���ݻ����uH�s H��H���J����H�� [^_]A\�H��薻��L�`L���L M��H��H������H�C ��H��H���{ H������H���N H�K H9�t
H��t�8L �3U H���P �Ɛ��������VSH��(1�H��H�A    H�����AH�R H��5 1�H��H�C �����H��([^�H��H���� H���L��������������SH�� H���   H��H�� [�K ������VSH��(H��Q H�q H�H���� H9�tH��tH���rK H�KH��tH��PH�K�J H��H��([^�l ������������VSH��(H�CQ H�q H�H���d H9�tH��tH���K H�KH��tH��PH�K�� H��H��([^� ������������VSH��8H��� H��H�L�D$/H��H�I�����H��8[^�H��H���h� H��� ������������������VSH��(H�c� H��H�L�BH��H�H�I��  �H��([^�H��H���� H��������������������H�� H��H�H��H�����������VSH��(H�CP H��H�H�I�����H�ı      ([^�H��H���� H���i�����������SH�� H���   H��H�� [��I ������SH��0H��O H�H��H�I�������A���~H���T� �H��0[�H�T$/H������H���7� �H��0[�SH�� H��H��H�I�{���H��H�� [Ð�SH�� H���#" H�,� H��H�H�� [Ð��������������SH�� H���C" H��� H��H�H�� [Ð��������������SH�� H���" H�<O H�H�� [Ð��SH�� H�$O H��H��" H��H�� [�H ������������H��N H��" �ATUWVSH��0��$�   L��D��H�L$ H�T$(��   H��vFL�d$ 1��   �@ =��  HF�H�{H��H9�s*��L���`  9�s�H�D$ H��0[^_]A\û   �    H9�u�H�L$ ����  ���  C����!  H�D$ H��0[^_]A\ÐL�d$ L���  �f�����������������SH�� �I��uH�� [�H��� �  ��tA�#�H�� [� H��� �  ��t�A��ǐ���������1�L�H�QL)�H��w��f� fA� �]� A�@�   H�Ð�������������   ��t+L�	1�L�AM)ȃ�t%I��v�� fA��   H��f.�     I��v��� fA��   H�Ð����VS�����L�L�IM)�tQE�E��yTA��������v=A���wSI�������t,E�H��E��A���A���uA��C��
����9�wI��L�[^�f�     I��A��L�[^�f�A���wjI�������v�E�H��E��A���A���u�A���uA���v�E�X�����D�ۃ�����u�A�      ��A��E�C������9�r�I��L��z���fD  A����j���I��������[���E�H��E��A���A����B���A���u
A����2���A���uA������������E�X�����D�ۃ���������A�X�ރ��@��������A��A��E�A��C�����7�9������I��L�������������������������L�L�IM)�I��vHA�A��fA��A��AD���D�� (��A���  v$D�� $��A���  vUA�   9�wK�BH��f�I��vJE�JE��fA��E��ED�E��E�� $��A���  w��
A�   A�� $��뱸�����f�     �����Ð�����������wH�H;A��   L�@L���   Á��  w<L�	1�L�AM)�I��v�I�AH�������@A�H���?�L�@L���   Á���  vc1����� w�L�	L�AM)�I��v�I�AH�������A�L�I�@H�������?���A� L�I�@H�������?���A� �D  L�	1�L�AM)�I���:���I�AH������� A��fD  1�Ð������������WVSH�� D��H��H��D�L$XH�T$X�q�������  ���  C�H�AH+H��vVH�H9Fu&�[9�r4H�H�JH�f�H�CH+H��v-H9Nt7D�D$X��H���������uȸ   H�� [^_�fD  1�H�� [^_�fD  �   H�� [^_Ð��WVSH�� A��H��H��D��uZH�H9CtaH�H9Fu'�4fD  9�r\H�H�JH��H�CH9t7H9Nt��H���w������uҸ   H�� [^_�D  �[   �f�     1�H�� [^_�fD  �      �   H�� [^_Ð��1�L�	L�AM)�I��v
E�fD9t� I���   L�	Ð��1�L�H�QL)�H��v��� fA9 t1����� A8@u�I���   L�Ð���SL�L9Y��   H�L�RI)�I����   E�A�� (��E�ځ��  vxE9�A��A��E��t1�ffD  L�RI)�I��vcE�[A�� (��E�ځ��  v<E9�w7E��fA��E��ED�fD�H�L�H��M�SL9QH�L�u�1�[�fD  �   [�f�     �   [Ð��������AUATUWVSH��(A��H��H��D����   A��D��L�.L�fM9�tXH�CH9tO��H�����������   9���   =��  H�H�Kw<H9�t@L�.��L�ff����D�H�JM9�H�f�u�1�H��([^_]A\A]��    H)�H��w�   L�.L�fH��([^_]A\A]É�f%���
f- $f��@(��uf��f��f�
H�JH�f�B�3���������"��� ��$�   1�������H��([^_]A\A]�f��   H��([^_]A\A]Ð�������������WVSH��0�D$pD��H�L$ H�T$(uUI�X�����  ���  C�M��t+H�|$ f�     ��H���f���9���H����H����u�H�D$ H��0[^_�fD  H�|$ L�D$`H���.���L�D$`뒐������UWVSH��(H��D��H��D�L$hH�T$h��������  ���  C�H��H�]�t+f�     D�D$h��H������9���H����H����u�H�H��([^_]Ð�H��8D�\$`A��I��t H��D�D$,H�T$ �����H�T$ ��D�D$,tE��L��H��8�   �   H��8Ð����WVSH�� H�I��H��D��D���W�      �     ����   H����   �@�� $�����  wi��
A�   �� $��9�wUH���o�����tkI�J�PI�M�CL��H)�H��H��I9�t<�D�� (��A���  v��� $��=�  v
9�A�   v��   H�� [^_�D  1�H�� [^_�fD  �   H�� [^_Ð��H��(H�	�ĭ���H��(�H��H��t����;@ �����������H�Ð�����������SH�� H��D��I����	��H��tH�; t1�H�� [�f.�     H��L�����H��H�t�H���CH�� [�H�	�Ь����������SH�� H��H�	H��t@�{ uH��H�    H�� [�f.�     蛬��H�    ��uH��H�� [��    1�H�� [Ð�������ATUWVSH�� L�%�4 H��H��D���@ A�ԃ8uH�������A��H�����k���Hc�H���t�H��H�� [^_]A\Ð�����������VSH��(H��L������I��H�ډ�H��([^��	��������������VSH��(H��D���_���A��H�ډ�����H��([^�H��H��t����> �������UWVSH��(H�9 H��H��uPH��tKH�5�3 �֋(���     �	f��փ8u)H���Y�����u��։(H��H��G H��([^_]�fD  �։(1�H��([^_]ÐVSH��(H��D��������H��tH�; t1�H��H��([^�fD  H���n���H��H�t܅��Cu�E1�A�   1�H���������H��H��t�#���= ��������������UWVSH��(L��H��H��L���'���H��u"L�D$pH����c��H�H��([^_]��    I��H�����C��H9�u�H�����������VSH��h1�H��������      H�T$ ����2 ��u�D$&f% �f= �tH��H��h[^�fD  H�\$8H������A�   1҉�����H)�H��H��h[^Ð������H�    �A Ð�������������������SH��0H�L�D$/H��H�1�1�购��H�H��0[Ð����������H��8L�L$/�����H��8Ð�����������L�BH�����������������������������������������SH��01�L�D$/H��1��:���H�H��0[ÐH��8�����H�	��A���~H��8�fD  H�T$/H�������H��8Ð�����������SH�� H������H��H�� [Ð���������SH�� H��賸��H��H�� [Ð���������H�AH�L�H�BI9�t-L�L�BL�AL�BL�AH�H�B    �B �f.�     �oBA�Ӑ����E1�H�AI�H��.	 ��������������E1�H�AH�H�L�BH��I���	 ����E1�H�AH�H�L�BH��I��	 ����H�L�B���������H�AH�A    H��A Ð�����������H�H�AH9�tH���7 Ð����������SH�� L�IH��H��H�H�L�CL9�tbL9�t=H�H�KH��L�HH�HH�KH�Ht4H�L�KH�C    � H�� [�f�     H�H�SH�PH�SH�PL�L����D  H��H��H�D$0� H�H�D$0묐�����SH�� H��� H��H�� [Ð���������UWVSH��(H�=�~ H��M��1�E1�H��H����� H�$= �   H���� ��tH�=�~ �   H����� ��u	H��([^_]�H�sH���B� E1�H��H����� �H��([^_]�H��H���� H������      ��������H��X�����������H��H�����������SH�� H��< H��H��9� H��H�� [��5 ������������H�Y< H��� �UWVSH��(H�=�} H��L��H���#� H��< �   H��H���� ��tH�=�} �   H����� ��uH��([^_]� H�sH���D� E1�H��H����� H��H��([^_]��� H��H��H��P H��� H��� H��H�PH��+� H���������H��8�����������H��(�����������SH�� H�tP H��H�H�I�� H�n� H��H��H���� H��H�� [�4 ��SH�� H�4P H��H�H�I�u� H�.� H��H��H�H�� [�� ����������SH�� H���s���H�L� H��H�H�� [Ð��������������SH�� H������H�� H��H�H�� [Ð��������������SH�� H�������H�\; H�H�� [Ð��SH�� H�D; H��H��	���H��H�� [��3 ������������H�; H�������SH�� H������H��� H��H�H�� [Ð��������������SH�� H�������H�l� H��H�H�� [Ð��������������SH�� H������H��: H�H�� [Ð��SH�� H��: H��H��I���H��H�� [�3 ������������H��: H��!����SH�� H�������H��� H��H�H�� [Ð��������������SH�� H������H��� H��H�H�� [Ð��������������SH�� H���S���H�<: H�H�� [Ð��SH�� H�$: H��H�����H��H�� [�L2 �������������      H��9 H��a����SH�� H�: H��H��	 H��H�� [�2 ������������H��9 H��� �SH��`H��$�   �Ao	H�ˋ�$�   L��L��t L�L�P)L$PH���d��L�L$@Ic�L�T$HL���f�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[�SH��`H��$�   �Ao	H�ˋ�$�   L��L��z L�L�P)L$PH���d��L�L$@Ic�L�T$HL���f�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[�SH��`H��$�   �Ao	H�ˋ�$�   L��L�.r L�L�P)L$PH���d��L�L$@Ic�L�T$HL���f�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H�      ��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[�SH��`H��$�   �Ao	H�ˋ�$�   L��L��w L�L�P)L$PH���d��L�L$@Ic�L�T$HL���f�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P(H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P8H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���P0H��H��`[�H��$�   L�L$@L�D$PH�L$0H��$�   H�L$(H��$�   H�L$ H���PH��H��`[�AWAVAUATUWVSH��   )�$�   H��$   I�)I�yL��$  �o8H��L��H��$   D��$  H��t_M�H�D$8L�L$PH��H��$  H�l$`L�D$`H�|$h)|$PL�d$0H�D$(D�|$ A�R�(�$�   H��H�Ę   [^_]A\A]A^A_�L�t$w1�1�L�l$xM���	���H�L$`H�l$PH��$  H�D$xH�L�L$@H�|$XL�D$P)|$@H�T$(H��L�l$8L�d$0D�|$ �PH�    �����D$hH!�H�l$`H	�A�$��t0H�L$xH�+�����H�{��A����D���H��L��膢���3�����      H��$(  H�@ H��t
H��$(  ��H��$(  L��襶��H�L$xH��$(  H�A�H�BH��H��  H�P �H��H�D$xL��H�H��,���H���T�������ATUWVSH��   H��$�   I�9I�YH��$�   �oL��H��H��$   L��$�   D��$�   L�H��tBL�L$(L�L$PD�D$ L�D$`H�|$`H�\$h)L$PH�D$8H�l$0A�RH��H�Đ   [^_]A\�L�d$pL�L$(I�D$D�D$ H�D$pH�L$`H�D$x    L�L$@Ƅ$�    L�D$PH�|$PH�\$X)L$@L�d$8H�l$0A�RH�    �����D$hH!�H�|$`H	ËE ��t)H�L$pI��H�>H�^L9��`����( �V���fD  H��$  H�@ H��t
H��$  ��H��$  E1�H��$  H�T$pL�D$xH��H�I��)� H��$  H�*  H�H �x���H�L$pI��H��L9�t�;( H���������AUATUWVSH��   )�$�   )�$�   H��$  �AoH��$(  ��$  �o8H��L��)D$@H��$0  H��t]M�H�D$8L�L$`H��H��$   )D$pL�D$p)|$`H�|$0�l$ H�D$(A�R�(�$�   H��(�$�   H�ĸ   [^_]A\A]�L��$�   1�1�L��$�   M������foT$@H�L$p)|$PH��$   L�l$8L�L$PH��$�   H�L�D$`)T$`H�|$0H�T$(H��l$ �PH�D$pH�D$@�fot$@f�t$x��t7H��$�   3�������A����<���H��L�������+���f�     H��$8  H�@ H��t
H��$8  ��H��$8  L���U0��H��$�   H��$8  H�A�H�BH��H�c  H�P �{���H��H��$�   L��H�H�      ���H�����������������WVSH��   )�$�   H��$�   �AoH��$  L��$   �oL��H��)D$@H��$  D��$�   L�H��tIL�L$(L�L$`D�D$ L�D$p)D$p)L$`H�D$8H�t$0A�R�(�$�   H��H�İ   [^_�fD  H��$�   fo\$@1�L�L$(H�Gf��$�   D�D$ H�L$pH��$�   L�L$P)\$`L�D$`HǄ$�       )L$PH�|$8H�t$0A�RH�D$pH�D$@�fot$@f�t$x��t"H��$�   H��3H9��N����% �D���H��$  H�@ H��t
H��$  ��H��$  E1�H��$  H��$�   H��H�H��$�   H��L�B� H��$  H�5�  H�p �u���H��$�   H��H��H9�t�~$ H�������������AUATUWVSH��   )|$pH��$�   �Ao9��$�   ��$�   �(H��L��H��$   H����   ��H�x  ��   L�@L�l$h��H�L�d$gL��M���,���H�)|$PH��H��$�   L�l$0D�͉\$(L�D$PH�T$ H���PH�L$h�������A���~Y(|$pH��H�Ĉ   [^_]A\A]ÐH�T$@I� ��)|$PH�T$0H��$�   D���|$@L�D$P�\$(H�T$ H���P�D  H��L��脛���H�[f ��� H��H�D$hL��H�H��r���H����������������ATUWVSH��   )�$�   H��$�   �Ao9D��$�   ��$�   �(H��L��H��$   H����   ��H�x  ��   H�H�t$`E1���L�@H�NH�L$`H��I��� �\$(H�E��)|$PL�D$PH��H��H��$�   H�t$0H�\$ �PH�L$`H��H9�t�`" �      �(�$�   H��H�Đ   [^_]A\�fD  I� H�T$@��)|$PH��$�   H�T$0E��H���|$@L�D$P�\$(H�t$ �P�H�.l �y� H�L$`H��H��H9�t��! H���K��������������AUATUWVSH��   )|$pH��$�   �Ao9��$�   ��$�   �(H��L��H��$   H����   ��H�x  ��   L�@L�l$h��H�L�d$gL��M���*��H�)|$PH��H��$�   L�l$0D�͉\$(L�D$PH�T$ H���PH�L$h�������A���~Y(|$pH��H�Ĉ   [^_]A\A]ÐH�T$@I� ��)|$PH�T$0H��$�   D���|$@L�D$P�\$(H�T$ H���P�D  H��L�������H��c �&� H��H�D$hL��H�H�����H�����������������ATUWVSH��   )�$�   H��$�   �Ao9D��$�   ��$�   �(H��L��H��$   H����   ��H�x  ��   H�HH�t$`E1���H�H�FH�D$`L�JH���R �\$(H�E��)|$PL�D$PH��H��H��$�   H�t$0H�\$ �PH�L$`H��H9�t� �(�$�   H��H�Đ   [^_]A\�D  I� H�T$@��)|$PH��$�   H�T$0E��H���|$@L�D$P�\$(H�t$ �P�H��i ��� H�L$`H��H��H9�t�C H�����������������SH�� H�� H��H�H�I��iuH��PH�� H�KH��H���� H����� H��H�� [�� �SH�� H�t H��H�H�I��iuH��PH�v� H�KH��H��� H���� H��H�� [� �SH�� H�� H��H�H�I��iuH��PH�f��       H�KH��H��6� H��H�� [�Y� ���������SH�� H�� H��H�H�I��iuH��PH�֮ H�KH��H���� H��H�� [�	� ���������SH�� H�� H��H�H�I��iuH��PH�ֱ H�KH��H��� H���� H��H�� [� �SH�� H�� H��H�H�I��iuH��PH�F� H�KH��H��F� H���n� H��H�� [�Q �SH�� H�$ H��H�H�I��iuH��PH�6� H�KH��H���� H��H�� [�� ���������SH�� H� H��H�H�I��iuH��PH��� H�KH��H��� H��H�� [��� ���������SH�� H� H��H�H�I ��iuH��PH���u� H��H�� [�x ��������SH�� H� H��H�H�I ��iuH��PH����c H��H�� [�8 ��������SH�� H�� H��H�H�I ��iuH��PH��H�� [�� SH�� H�� H��H�H�I ��iuH��PH��H�� [�pc SH�� H�� H��H�H�I ��iuH��PH���e� H��H�� [� ��������SH�� H�� H��H�H�I ��iuH��PH����d H��H�� [�X ��������SH�� H�$ H��H�H�I ��iuH��PH��H�� [��� SH�� H�4 H��H�H�I ��iuH��PH��H�� [�`d SH�� H�D H�H�A H��H�@    H�I��iuH��PH���� H��H�� [� ������������SH�� H�D H�H�A H��H�@    H�I��iuH��PH�      ���Ig H��H�� [�\ ������������SH�� H�� H�H�A H��H�@    H�I��iuH��PH��H�� [�D� ����SH�� H�� H�H�A H��H�@    H�I��iuH��PH��H�� [�f ����SH�� H�� H�H�A H��H�IH�@    ��iuH��PH���9� H��H�� [� ������������SH�� H�� H�H�A H��H�IH�@    ��iuH��PH���i H��H�� [�< ������������SH�� H�$ H�H�A H��H�IH�@    ��iuH��PH��H�� [锚 ����SH�� H�4 H�H�A H��H�IH�@    ��iuH��PH��H�� [�i ����SH�� H�D H��H�H�I��iuH��PH�� H��H��H��� H��H�� [�j ����������SH�� H�D H��H�H�I��iuH��PH�6� H��H��H��7� H��H�� [� ����������SH�� H��
 H��H�H�I��iuH��PH�v� H��H��H�H�� [��� ��SH�� H��
 H��H�H�I��iuH��PH��� H��H��H�H�� [�� ��SH�� H��
 H��H�H�I��iuH��PH�� H��H��H��g� H��H�� [�J ����������SH�� H��
 H��H�H�I��iuH��PH�&� H��H��H��� H��H�� [�� ����������SH�� H�4
 H��H�H�I��iuH��PH�f� H��H��H�H�� [��� ��SH�� H�D
 H��H�H�I��iuH��PH��� H��H��H�H�� �      [�� ��SH�� H�d
 H��H�H�I��iuH��PH�F� H��H��H��G� H��H�� [�* ����������SH�� H�D
 H��H�H�I��iuH��PH�� H��H��H���� H��H�� [�� ����������SH�� H��	 H��H�H�I��iuH��PH��� H��H��H�H�� [�� ��SH�� H��	 H��H�H�I��iuH��PH��� H��H��H�H�� [�b� ��SH�� H��	 H��H�H�I��iuH��PH�6� H��H��H��'� H��H�� [�
 ����������SH�� H��	 H��H�H�I��iuH��PH�� H��H��H���� H��H�� [� ����������SH�� H�	 H��H�H�I��iuH��PH��� H��H��H�H�� [�� ��SH�� H�� H��H�H�I��iuH��PH�v� H��H��H�H�� [�B� ��SH�� H�� H��H�H�I��iuH��PH�&� H��H��H��� H��H�� [�� ����������SH�� H�� H��H�H�I��iuH��PH��� H��H��H��� H��H�� [� ����������SH�� H�D H��H�H�I��iuH��PH��� H��H��H�H�� [�b� ��SH�� H�4 H��H�H�I��iuH��PH�f� H��H��H�H�� [�"� ��SH�� H�$ H��H�H�I��iuH��PH�� H��H��H���� H��H�� [�� ����������SH�� H� H��H�H�I��iuH��PH�� H��H��H��� H��H�� �      [�z ����������SH�� H�� H��H�H�I��iuH��PH�v� H��H��H�H�� [�B� ��SH�� H�t H��H�H�I��iuH��PH�V� H��H��H�H�� [�� ��SH�� H�d H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH������H��H�� [� ��������SH�� H�d H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH���e� H��H�� [� ��������SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [�0���SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [�� SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH���5���H��H�� [�� ��������SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH���� H��H�� [�x ��������SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [�P���SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [�� SH�� H�� H�H�A H��H�@    H�A H�@0  �        H�A H�@@    H�A H�@P    H�I��iuH��PH���e���H��H�� [�H ��������SH�� H�� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH���� H��H�� [�� ��������SH�� H� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [逭��SH�� H� H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [��� SH�� H�$ H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��蕰��H��H�� [� ��������SH�� H�$ H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH����� H��H�� [�8 ��������SH�� H�D H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [鰯��SH�� H�T H�H�A H��H�@    H�A H�@0    H�A H�@@    H�A H�@P    H�I��iuH��PH��H�� [�� H��8�����H�	��A���~H��8�fD  H�T$/H���r����H��8Ð�����������H�H�AH9�tH��� Ð����������H��8�����H�	��A���~H��8�fD  H�T$/H�������H��8Ð�����������H�H�AH9�tH���
 Ð����������ATUWVSH��PH��L��H��$�   E��L��$��         H�l$@L�L$>H��H�t$H視��H�H�l$(E����$�   H��D��$�   �T$ H���PH�C H��tH����H��H��趖��H�L$HH�A�H�CH�����H�C �������A���~ H�L$@�������A���~H��P[^_]A\�f�H�T$?H��������H��H�������H��P[^_]A\�H�T$?H��H�D$HH�H�����H�D$@H��H�H�����H���	���H���␐��ATUWVSH��pH��L��H��$�   E��L��$�   H�\$0E1�H�CH��H�D$0H�|$PI��L� H�E E��H����$�   H�\$(D��$�   �T$ H���PH�F H��tH����H�T$PH�FE1�H��L�D$XH�I��� H�L$PH�����H��H�F H9�t�� H�L$0H��H9�t�� �H��p[^_]A\�H��H�L$0H��H9�t� H������H�L$PH��H��H9�t�� �͐���ATUWVSH��PH��L��H��$�   E��L��$�   H�l$@L�L$>H��H�t$H���H�H�l$(E����$�   H��D��$�   �T$ H���PH�C H��tH����H��H������H�L$HH�A�H�CH�����H�C �������A���~ H�L$@�������A���~H��P[^_]A\�f�H�T$?H���������H��H��������H��P[^_]A\�H�T$?H��H�D$HH�H�����H�D$@H��H�H�����H�������H���␐��ATUWVSH��pH�\$0H��H��$�   E��H�CE1�H��H�D$0H��$�   L��H�|$PL�B�k  H�E E��H����$�   H�\$(D��$�   �T$ H���PH�F H��tH����H�FH�T$PE1�H��H�H�D$XL�B��  H�L$PH�����H��H�F H9�t� H�L$0H��H9�t��      � �H��p[^_]A\�H��H�L$0H��H9�t�r H�������H�L$PH��H��H9�t��T �͐�WVSH��@H�t$8H��L��H�|$7M��H��I���[���H�H��H��L��$�   �PH�L$8�������Q���~H��@[^_�H��H���D$,�~���D$,H��@[^_�H��H�D$8H��H�H��~��H���4�������VSH��XH�\$0H��L��H�CH��O�E1�H�D$0�� H�H��H��L��$�   �PH�L$0H��H9�t�D$,�l �D$,H��X[^�H�L$0H��H��H9�t�K H���������WVSH��@H�t$8H��L��H�|$7M��H��I���K���H�H��H��L��$�   �PH�L$8�������Q���~H��@[^_�H��H���D$,�}���D$,H��@[^_�H��H�D$8H��H�H���|��H���$�������VSH��XH�\$0H��L��H�CH��O�E1�H�D$0�� H�H��H��L��$�   �PH�L$0H��H9�t�D$,�\ �D$,H��X[^�H�L$0H��H��H9�t�; H���������H�H�@ H��D��H��H�H�@ H��D��H��H�H�@ H��D��H��H�H�@ H��D��H��L�T$0H��L��M��L�L$(H�L�T$(H�`�L�T$0H��L��M��L�L$(H�L�T$(H�`�L�T$0H��L��M��L�L$(H�L�T$(H�`�L�T$0H��L��M��L�L$(H�L�T$(H�`�VSH��8H�H�t$(L��M��L�L$pH���PH�C H��tH����H��H��踏��H�L$(H�A�H�CH�����H�C �������A���~H��8[^�H�T$'H���-{���H��8[^�H�T$'H��H�D$(H�H��{��H���G����������VSH��HH�H�t$ L��M��L��$�   H���PH�C H��tH�����      H�T$ H�CE1�H��L�D$(H�I��A� H�L$ H�E���H��H�C H9�t�c �H��H[^�H�L$ H��H��H9�t�E H�������������������VSH��8H�H�t$(L��M��L�L$pH���PH�C H��tH����H��H�����H�L$(H�A�H�CH�����H�C �������A���~H��8[^�H�T$'H��������H��8[^�H�T$'H��H�D$(H�H������H�������������VSH��HH�H�t$ L��M��L��$�   H���PH�C H��tH����H�CH�T$ E1�H��H�H�D$(L�B�@� H�L$ H�d���H��H�C H9�t�" �H��H[^�H�L$ H��H��H9�t� H���l���������������H�H�@H��H�����H�H�@H��H�����H�H�@H��H�����H�H�@H��H�����ATUWVSH��0H�L��H��H���PH�|$(H��CHH��Pƃ�   H��H��CIH�C    H�C(    H�C8    H��P H�D$(H�h�H�M�f  E1�I��H��H��I������H�L$(A�, �����L�cH�k��A�����   H�H��H���P(H�D$(H�h�H�M�  E1�I��H��H��I���|��H�L$(A�, �����L�c(H�k0��A�����   H�H��H���P0H�D$(H�p�H�N�� E1�I��H��H��H���&��H�L$(�D5  �����H�k8H�s@��A���~&H��0[^_]A\�H�T$'H���}w���:����     H�T$'H���bw���H��0[^_]A\�fD  H�T$'H���Bw���U���H�T$'H��H�D$(H�H��7w��H���_������ސ����������ATUWVSH��@H�L��H��H���PH�t$ H���CHH��Pƃ�   H��H����      CIH�C    H�C(    H�C8    H��P H�l$(H�M�� E1�I��H��H��I���6���H�L$ H�FA�, L�cH�kH9�t�F� H�H��H���P(H�l$(H�M�L� E1�I��H��H��I������H�L$ H�FA�, L�c(H�k0H9�t��� H�H��H���P0H�|$(H�O��� E1�I��H��H��H��蚘��H�L$ H���D=  H�k8H�{@H9�t�� �H��@[^_]A\�H�L$ H��H��H9�t�� H����������ސ�����������AUATUWVSH��8H�L��H��H���PH�|$(H��f�CHH��PH��ƃ�   H��f�CJH�H�C    H�C(    H�C8    �P H�D$(H�h�H�M�"� E1�I��H��H��I�����H�L$(A�, �����L�cH�k��A�����   H�H��H���P(H�D$(L�`�H��������?I�L$H9��J  H�,	H���� E1�M��H��H��I�������H�L$(1�L�k(�����fA�T-�L�c0��A�����   H�H��H���P0H�D$(H�h�H��������?H�uH9���   H�H���?� E1�I��H��H��I���{���H�L$(1�L�c8fA�D4������H�k@��A���~;H��8[^_]A\A]�H�T$'H����s��������     H�T$'H��������W���H�T$'H�������H��8[^_]A\A]�H�T$'H��H�D$(H�H�����H�������H�T$'H��H�D$(H�H��s��H���������� �	 ���������AUATUWVSH��HH�L��H��H���PH�t$ H��f�CHH��PH��ƃ�   H��f�CJH�H�C    H�C(    H�C8    �P H�l$(H�M��� E1�I��H��H��I��蒕��H�L$ H�FA�, L�c�      H�kH9�t�� H�H��H���P(L�d$(H��������?I�L$H9���   H�,	H���� E1�M��H��H��I��艢��H�L$ H�F1�L�k(fA�T-�L�c0H9�t�6� H�H��H���P0H�l$(H��������?H�}H9�wwH�H���'� E1�I��H��H��I���#���H�L$ H��1�L�c8fA�D<�H�k@H9�t��� �H��H[^_]A\A]�H�L$ H��H��H9�t�� H�����������[ �V ������ATUWVSH��0H�L��H��H���PH�|$(H��C!H��PH��C"H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CoH��P H�D$(H�h�H�M�5� E1�I��H��H��I�����H�L$(A�, �����L�cH�k��A����!  H�H��H���P(H�D$(H�h�H�M��� E1�I��H��H��I���K��H�L$(A�, �����L�c(H�k0��A����
  H�H��H���P0H�D$(H�h�H�M�� E1�I��H��H��I���� ��H�L$(A�, �����L�c8H�k@��A�����   H�H��H���P8H�D$(H�h�H�M�3� E1�I��H��H��I��� ��H�L$(A�, �����L�cHH�kP��A���~?H�H���PHH��C\H��PP�C`H��0[^_]A\�H�T$'H����o�������f�     H�T$'H����o���H�T$'H���o���L���H�T$'H���o�������H�T$'H��H�D$(H�H��o��H��輾�������ܐ�����ATUWVSH��@H�L��H��H���PH�|$ H��C!H��PH��C"H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CoH��P H�l$(H�M��� E1�I��H��H��I����      ���H�L$ H�GA�, L�cH�kH9�t�� H�H��H���P(H�l$(H�M�� E1�I��H��H��I���7���H�L$ H�GA�, L�c(H�k0H9�t�G� H�H��H���P0H�l$(H�M�M� E1�I��H��H��I������H�L$ H�GA�, L�c8H�k@H9�t��� H�H��H���P8H�l$(H�M��� E1�I��H��H��I��蛐��H�L$ H��A�, L�cHH�kPH9�t�� H�H���PHH��C\H��PP�C`H��@[^_]A\�H�L$ H��H��H9�t�r� H���ڼ�������ܐ���ATUWVSH��0H�L��H��H���PH�|$(H��C!H��PH��C"H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CoH��P H�D$(H�h�H�M�� E1�I��H��H��I���q���H�L$(A�, �����L�cH�k��A����!  H�H��H���P(H�D$(H�h�H�M�� E1�I��H��H��I������H�L$(A�, �����L�c(H�k0��A����
  H�H��H���P0H�D$(H�h�H�M�Y� E1�I��H��H��I�������H�L$(A�, �����L�c8H�k@��A�����   H�H��H���P8H�D$(H�h�H�M�� E1�I��H��H��I���o���H�L$(A�, �����L�cHH�kP��A���~?H�H���PHH��C\H��PP�C`H��0[^_]A\�H�T$'H���k�������f�     H�T$'H���k���H�T$'H���k���L���H�T$'H���ok�������H�T$'H��H�D$(H�H��dk��H��茺�������ܐ�����ATUWVSH��@H�L��H��H���PH�|$ H��C!H��PH��C"H��P@H�C    H��H��CXH�C(    H�      �C8    H�CH    �CoH��P H�l$(H�M�� E1�I��H��H��I���U���H�L$ H�GA�, L�cH�kH9�t�e� H�H��H���P(H�l$(H�M�k� E1�I��H��H��I������H�L$ H�GA�, L�c(H�k0H9�t�� H�H��H���P0H�l$(H�M�� E1�I��H��H��I��蹌��H�L$ H�GA�, L�c8H�k@H9�t��� H�H��H���P8H�l$(H�M��� E1�I��H��H��I���k���H�L$ H��A�, L�cHH�kPH9�t�{� H�H���PHH��C\H��PP�C`H��@[^_]A\�H�L$ H��H��H9�t�B� H��誸�������ܐ���AUATUWVSH��8H�L��H��H���PH�|$(H��f�C"H��PH��f�C$H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CzH��P H�D$(H�h�H�M��� E1�I��H��H��I���=���H�L$(A�, �����L�cH�k��A����|  H�H��H���P(H�D$(L�`�H��������?I�L$H9���  H�,	H���`� E1�M��H��H��I������1�L�k(�����fA�L-�H�L$(L�c0��A����%  H�H��H���P0H�D$(L�`�H��������?I�l$H9��|  H�H����� E1�M��H��H��I���)���H�L$(1�L�k8�����fA�T-�L�c@��A�����   H�H��H���P8H�D$(L�`�H��������?I�L$H9��  H�,	H���y� E1�M��H��H��I������H�L$(1�L�kHfA�D-������L�cP��A���~rH�H���PHH��C\H��PP�C`H��8[^_]A\A]�H�T$'H���g���q���f.�     H�T$'H������������H�T$'�      H��������(���f.�     H�T$'H��������{���H�T$'H��H�D$(H�H���f��H������H�T$'H��H�D$(H�H�����H���ѵ���� �� ������ ��������������AUATUWVSH��HH�L��H��H���PH�|$ H��f�C"H��PH��f�C$H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CzH��P H�l$(H�M��� E1�I��H��H��I��聈��H�L$ H�GA�, L�cH�kH9�t�� H�H��H���P(L�d$(H��������?I�L$H9��m  H�,	H���|� E1�M��H��H��I���x���H�G1�L�k(fA�L-�H�L$ L�c0H9�t�%� H�H��H���P0L�d$(H��������?I�l$H9���   H�H���� E1�M��H��H��I������H�L$ H�G1�L�k8fA�T-�L�c@H9�t�� H�H��H���P8L�d$(H��������?I�L$H9���   H�,	H���� E1�M��H��H��I��衔��H�L$ H��1�L�kHfA�D-�L�cPH9�t�N� H�H���PHH��C\H��PP�C`H��H[^_]A\A]�H�L$ H��H��H9�t�� H���{�������� ���� ���� ������AUATUWVSH��8H�L��H��H���PH�|$(H��f�C"H��PH��f�C$H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CzH��P H�D$(H�h�H�M�� E1�I��H��H��I�������H�L$(A�, �����L�cH�k��A����|  H�H��H���P(H�D$(L�`�H��������?I�L$H9���  H�,	H��� � E1�M��H��H��I���\���1�L�k(�����fA�L-�H�L$(L�c0��      �A����%  H�H��H���P0H�D$(L�`�H��������?I�l$H9��|  H�H���� E1�M��H��H��I�������H�L$(1�L�k8�����fA�T-�L�c@��A�����   H�H��H���P8H�D$(L�`�H��������?I�L$H9��  H�,	H���9� E1�M��H��H��I���u���H�L$(1�L�kHfA�D-������L�cP��A���~rH�H���PHH��C\H��PP�C`H��8[^_]A\A]�H�T$'H����a���q���f.�     H�T$'H�����������H�T$'H�������(���f.�     H�T$'H�������{���H�T$'H��H�D$(H�H��a��H��诰��H�T$'H��H�D$(H�H��Y���H��葰����� ��� ������� ��������������AUATUWVSH��HH�L��H��H���PH�|$ H��f�C"H��PH��f�C$H��P@H�C    H��H��CXH�C(    H�C8    H�CH    �CzH��P H�l$(H�M�� E1�I��H��H��I���A���H�L$ H�GA�, L�cH�kH9�t�Q� H�H��H���P(L�d$(H��������?I�L$H9��m  H�,	H���<� E1�M��H��H��I���8���H�G1�L�k(fA�L-�H�L$ L�c0H9�t��� H�H��H���P0L�d$(H��������?I�l$H9���   H�H����� E1�M��H��H��I���͏��H�L$ H�G1�L�k8fA�T-�L�c@H9�t�z� H�H��H���P8L�d$(H��������?I�L$H9���   H�,	H���e� E1�M��H��H��I���a���H�L$ H��1�L�kHfA�D-�L�cPH9�t�� H�H���PHH��C\H��PP�C`H��H[^_]A\A]�H�L$ H��H��H9�t�      ��� H���;������� ���}� ���v� ������SH�� H��� H��H�H�I 赚 H��� H��H�胴��H��H�� [�v� ������SH�� H��� H��H�H�I �u� H��� H��H�H�� [�>������������������   �6� ������Ð��������������D�AXH�AhA��H�AH�At*H��~%H�H�AH�A(    H�A     H�A0    �D  A��H�At�H��u�H�QpH��v�H�A(H�A H�D�H�A0Ð����VSH��8H��H���   H��H��P0��tH�C+CH��8[^�D  H���   H��H�CH+CL���   L�L���   H�D$ A�R8H�H��   +��   H��8[^Ð����������������    u1H�AƁ�   H���   H�AH���   H�A{H�AH�AH�A|H�AÐ�������    t:H�AƁ�    H9AH���   L�Ah����H��   H�QL�AH���   H�AÐ�����������AWAVAUATUWVSH���   �   H�A(H9A H��sH�������Ph���@�ƀ{z txH���   H����   H��P0��A��u[@��tVL�c`H�|$@H�l$8L�sHH���   L��$�   I��L��H�H�l$ �P����t��v3H������H���Ph���A��D���H���   [^_]A\A]A^A_�D  L�|$8I)�M��~�M��H��L��襧��I9�u��x�����0� ����������������UAWAVAUATWVSH��hH��$�   H��H���   H��L��H���.  H��P0��uqH���   H��P@Hc�H��H�BH���褦��H���   L�c`H)�H�I��L�t$@L�m�L�L�t$(L�}�H�T$0L��L�l$8L�7L�|$ �P���      v/����   H�KHI��H���Ŧ��H9���H�e�[^_A\A]A^A_]�L�U�H�{HL��E�H��L��L�U�L)�I��苦��H9�u�D�M�L�U�A��t�H���   L��L�K(L�E�H�L�l$8L�T$0L�t$(L�|$ �P��tH�u�L��H��L)�I���2����h���H�60 �1� 輍 ������������SH�� �yx H��tH�IhH��t��� H�Ch    �Cx H���   H��t��� Hǃ�       Hǃ�       Hǃ�       Hǃ�       H�� [Ð����SH�� �yx H��uH�yh tH�� [�D  H�Ip�� �CxH�Ch�␐�����������UWVSH��HH�qHH��H��H��D���������   A��  A��H��H������H���o������   �{x H�Chu	H����   H�C1�@��H�CH�C�C\�{Xf�SyH�C(    H�C     H�C0    �C`�Cdt#H�E1��|$ A�   H�L$0H���P H�|$0�tH��H��H[^_]�f�     H���x  1�H��H[^_]�H�Kp�� �CxH�Ch�c����������H��������������ATUWVSH��0H�AL�a8H��H�RH��H�|$(H�k8H�QH�SH�CH�AH�QH�SH�CH�AH�QH�S H�CH�A H�Q H�S(H�C H�A(H�Q(H�S0H�C(H�A0H�Q0L��H��H�C0�8� H��L���-� H��H���"� H���� H�FHH�SHH�VH�SPH�CH�FP�VP�SX�CP�FX�VX�S\�CX�F\�V\�S`�C\�F`�V`�Sd�C`�Fd�VdH�Sh�CdH�FhH�VhH�SpH�ChH�FpH�VpH�Cp�Fx�Sx�VxH���   �CxH���   H���   H���   H���   H���   H���   H���   H���   H���   �      H���   H���   H���   H���   H���   �SyH���   �Fy�Vy�Sz�Cy�Fz�VzH���   �CzH���   H���   H���   H���   H���   H���   ���   H���   ���   ���   ���   H��0[^_]A\Ð����H��(1�H�Q(H9Q sH�������Ph���������H��(Ð����WVSH��0H�yHH��H���J��������   H��H�\$(�S�������H�L$(�AX    Ɓ�    ����H�T$(1�H��f�ByH�BhH�B(    H�B     H�B0    H�BH�BH�B�B\�B`�Bd� ��H��t@��H��uH��0[^_�1�H��0[^_�H��H��u�� H��荠���8� �� �� �[���H���� H�L$(�W� H��菤��H���鐐��������WVSH��@H��H��H���� ���  H���{� H��H�KH�/������   �{y ��   H���   H����  H��P(�����   �{y ��   H���   H����  H��P0����   H��twH�H���P0��u&�SXE1�A�   H�H�L$0�T$ H���P H�|$0�tDH���   H��@[^_À{z �h���H���   H��@[^_�fD  �{z t�H����������   1�H���   H��@[^_�f�     1�����f�     H���   H�SdH���   H�CH+CL�I��L���   H�D$ A�R8Hc�H�H���   H���   H)���   H���   H�C(    H�C     H�C0    H�H���   H�ChH���   H�CH�CH�C�C\�C`�Cd�����D  H�ChH�C(    H�C     H�C0    H�CH�CH�C����� H���   I���iJ���i���藆 ��������      WVSH�� H��H��L��H�IH�'����uH��H	�uH�Cp   H��H�� [^_��     H��t�H��~�H��H�shH�{pH�� [^_Ð��ATUWVSH�� ���    H��H��L����   1�M��H�AH�Q~	H9���   H9�H�Khƃ�    ��H���   ��H��   D�cXH�KH�SH���   H�CH�{p�   HCCpH��H9�~$H���   H����  H��P0A��t����   I��H��H���e H�H��H�� [^_]A\�@ �yz uJD�aX1��f�� H�OH���H�CH�����    H�C�  D�cXH�Ͻ   �Z���f�     H�������Ph���t@H�Ch�Cz 1�D�cXH�C(    H�C     H�C0    H�CH�CH�C�
���f�     1��G���f�     H�SL�cI)�u8L�cH�H�H)�t!H�I��H��L��脜��H���t_H��u�H��u$�Cy�����H��M��L��-H��L�L)�Lc뮐H�ChH�C(    H�C     H�C0    �Cy H�CH�CH�C����H�X& 胅 �� H�SH�Ͻ   �����������������UWVSH��8�AXH��H���   H��L��@��H����   H��P0��t~@��ty�{y usL�C(H�C0L)��{z uH�SpH�J�H��HG�H=   �   HM�H9�>H�S H�t$ H�KHI��I)�L���"���H�H9�t:H��H)�H9Ÿ    HL�H��8[^_]�I��H��H��H��8[^_]�� f�     �KXH�Sh��H�SH�SH�Su��t!H�KpH��vH�S(H�S H�T
�H�S0�Cz�H�C(    H�C     H�C0    ���Â ���UWVSH��8H�����H��H��L���A    H��D���f��      ����uH��H��8[^_]�fD  H�NHA��H������H���t�1ҋ�$�   H�H��f�VyH���   H�F(    H�F     H�F0    H���   H���   H�Vh�~`�{H�VH�VH�VH��8[^_]Ð�����������AVAUATUWVSH��pH��H���   H��M��E��H����   H��    �P(��I�@��M��H�����L�sH���F    L��!��P ��<u@��tH��H��p[^_]A\A]A^�D  A��uzM��uu�{z tH���   H��P0��t^�C\1��{y �D$l��   �{z tH�{(H+{ 1�A�   L��轙��H���t�HǋD$lH�>�F��     �   1��B���@ ���    t:H�Cƃ�    H9CH���   H�Kh����H��   H�SH�KH���   H�CLcŋC\M�Ā{y �D$lu)�D$ H�L$PE��H�������H�D$PH��D$X�F������A��uыCdH�T$lH��L�D$8�D$l�!���L�D$8H�I��D$l먐�CdH�T$lH�ىD$l�����Hc����������UWVSH��HI�8I�hH�����H��H���A    H�JH������ti���    t:H�Cƃ�    H9CH���   H�Kh����H��   H�SH�KH���   H�CH�L$0�l$ E1�I��H�������H�D$0H��D$8�FH��H��H[^_]Ð����������VSH��X�AXH�ˉ���  �yy tx���    t:H�AH9AH���   ����H��   H���   H�IhH�CH�Sƃ�    H�KH�SdH��������SdH�L$0A�   Lc��T$ H���9���H�|$0��/  H�S L�C(L9�sp���tA�0H�C(H�S L�@L�C(I)�H����������   �SXH�Ch��H�CH�CH�C�      uN��uIH�C(    H�C     H�C0    �����t!H��X[^�f�H�SpH��w6���@�t$Ou|�Cz1�H��X[^�H�SpH��v�H�C(H�C H�D�H�C0�f��KXH�Ch��H�CH�CH�Cu��tcH�C(H�C H�D�H�C0����Czt�H�C(@�0��H�C(H��X[^�@ H�T$OA�   H��������t�Cz���E��������H��X[^�f�H�C(    H�C     H�C0    딐�����WVSH��@�AXH�ˉ��  �yz ��   H�AH;A���   ��   H�P�H�Q�P�1����tR9��tL@����   ���    H�Cu-H���   H�CH�S|H�Sƃ�   H���   H�C{H�CH�C�Cy@�0��H��@[^_�H�������Ph���trH�ChH�C(    ���   H�C     H�C0    �Cz H�CH�CH�CH�H�L$0H���D$    A�   I�������P H�|$0�tH�H���PH���������������l�����UWVSH��(�qX@��H��t|H�iHH���������tlH���   ��H�{H+{H��t^H��P(��x��uH��H��([^_]�H���#���H���   H��H��P@Hc�H��H�H��H�H��H��([^_]�f�     H���������{ ��AUATUWVSH��X�AXH���3  �yz �-  ���    H�A�e  H�SH9���  H���   �   H�{pHCspH��H�~���  H��P0���  H���   H��P(���i  Hc�H��H��H���   I��H���   H)�I)�H9�    LN�{y H���   tH�KH9K��  H9���  H��L���   ��  �C`M�4M��L���   L���   �Cd��  L�S1�M9�L�T$Hv�      o1�D  H���   L�D$HH�S`H�L�D$8M�:L�D$0L���   L�D$ M��L�T$(�P ������  L�L$HL+K��M����  M����	���(  L���   A�   L��H+��   L�H;��   �o  H�KHM��L������H����  H�����  1�H��   L���   L�SI��H���   L9�L�T$H�#������  @���y���H�Ch��H�C(    H�C     H�C0    �Cy H�CH�CH�C�  H�M ��z H�������Ph���t{H�ChH�C(    ���    H�C     H�C0    �Cz H�CH�CH�C�����H9Cƃ�    H���   H�Kh����H��   H�SH�KH9�H���   H�C�i���� H��X[^_]A\A]��     H���   H��P@H�H�l�H������@ L���   L�SH���   I)�L9�M��L��r0M��u1M��H���   �   ��	��2���f��   �y���fD  I��H��I��L���<��H���   H�� H�SH�KHI���0���H��I����   H�+ �y fD  M���  H�Ch�CXH�CH�C��   N� L�KH�C(    H�C     H�C0    �Cy� �����D  M���@��uH�O �y f.�     H�ChH�C(    H�C     H�C0    �Cy H�CH�CH�C���������f.�     H�C�n����    H����� H��I��urH���   H��t�� L���   H���   �D���1������H��tYH9�/L���   E1�I��L���:��L���   ����@��������+���H��E1��Q� I��H���   I��L���:���w���H9�~�H��      ��*� I���b���H�� �x �v �VSH��(H��H����  H�X� H�F@    H�H�CHH�FH�CP�FP�CXH�CH    �CP �CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �Fx�Cy�Cy �Fy�Cz�Cz �Fz�C{�F{H���   Hǃ�       H���   H���   Hǃ�       H���   ���   ƃ�    ���   H���   H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H�ChH�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��([^Ð����������ATUWVSH�� L�%�[ I�D$H�q8H��H�H�A    H�{HH�A    H�A    H�A     H�A(    H�A0    H���t� H�m� H��H�C@    H�H�S@����H�CX    H��H�C`    H�Ch    H�Cp   �Cx    Hǃ�       Hǃ�       ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       �C� ��uH�� [^_]A\�@ H���Ț H���   H�� [^_]A\�H��H���[���I�T$H��H��K� H���s������VSH��(H��H����  H�h� H�F@    H�H�CHH�FH�CP�FP�CXH�CH    �CP �CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �Fx�Cy�Cy �Fy�Cz�Cz �Fz�C{�F{H���   Hǃ�       H���   H���   Hǃ�       H���   ���   ƃ�    ����         H���   H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H�ChH�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��([^Ð����������ATUWVSH�� L�%�X I�D$H�q8H��H�H�A    H�{HH�A    H�A    H�A     H�A(    H�A0    H��脁 H�}� H��H�C@    H�H�S@����H�CX    H��H�C`    H�Ch    H�Cp   �Cx    Hǃ�       Hǃ�       ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       �S� ��uH�� [^_]A\�@ H���ؗ H���   H�� [^_]A\�H��H���k���I�T$H��H��[� H��背�����SH�� H��� H��H������H�KH�0���H��W H�K8H��H��� H��H�� [��� ������������SH�� H�4� H��H�����H�KH�����H�IW H�K8H��H�H�� [�Ā ����SH�� H��� H��H��Y���H�KH蠊��H�	W H�K8H��H�H�� [鄀 ����VSH��(H��H������H��H�����  H�SHH�FHH�VH�SPH�CH�FP�VP�CP�CX�CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �FxH���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   �Cy�Cy �Fy�Cz�Cz �FzH���   Hǃ�       H���   H���   H��      ��       H���   ���   ƃ�    ���   H�ChH�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��H��([^ÐD�AXH�AhA��H�AH�At*H��~%H�PH�AH�A(    H�A     H�A0    �@ A��H�At�H��u�H�QpH��v�H�A(H�A H�DP�H�A0Ð����VSH��8H��H���   H��H��P0��tH�CH+CH��H��8[^ÐH���   H��H�CH+CL���   L�L���   H��H�D$ A�R8H�H��   +��   H��8[^Ð�������������    u1H�AƁ�   H���   H�AH���   H�A|H�AH�AH�A~H�AÐ�������    t=H�A1�Ɓ�    H9AH���   L�Ah��H�PH���   H���   L�AH�AH�QÐ��������AWAVAUATUWVSH���   �   H�A(H9A H��sH����  �Phf���@�ƀ{z tyH���   H����   H��P0��A��u\@��tWL�c`H�|$@H�l$8L�sHH���   L��$�   I��L��H�H�l$ �P����t��v2H����  H���Phf���A��D���H���   [^_]A\A]A^A_� L�|$8I)�M��~�M��H��L���U���I9�uă��y������k ����������������UAWAVAUATWVSH��hH��$�   H��H���   H��L��H���.  H��P0��uqH���   H��P@Hc�H��H�BH����T���H���   L�c`H)�H�I��L�t$@L�m�L�L�t$(L�}�H�T$0L��L�l$8L�wL�|$ �P��v/����   H�KHI��H���u���H9���H�e�[^_A\A]A^A_]�L�U�H�{HL��E�H��L��L�U�L)�I���;���H9�u�D�M�L�U�A��t��      H���   L��L�K(L�E�H�L�l$8L�T$0L�t$(L�|$ �P��tH�u�L��H��L)�I�������h���H�� ��k �lj ������������SH�� �yx H��tH�IhH��t蔾 H�Ch    �Cx H���   H��t�w� Hǃ�       Hǃ�       Hǃ�       Hǃ�       H�� [Ð�����yx uH�yh t�f��   �����������SH�� H��������?H��H�IpH9�wH��-� �CxH�ChH�� [��� ����������UWVSH��HH�qHH��H��H��D���#�������   A��  A��H��H��藀��H�����������   �{x H�ChuH��uH���`���H�ChH�C1�@��H�CH�C�C\�{Xf�SyH�C(    H�C     H�C0    �C`�Cdt#H�E1��|$ A�   H�L$0H���P H�|$0�tH��H��H[^_]ÐH���h  1�H��H[^_]Ð������������H�������������ATUWVSH��0H�AL�a8H��H�RH��H�|$(H�k8H�QH�SH�CH�AH�QH�SH�CH�AH�QH�S H�CH�A H�Q H�S(H�C H�A(H�Q(H�S0H�C(H�A0H�Q0L��H��H�C0��w H��L����x H��H����x H���x H�FHH�SHH�VH�SPH�CH�FP�VP�SX�CP�FX�VX�S\�CX�F\�V\�S`�C\�F`�V`�Sd�C`�Fd�VdH�Sh�CdH�FhH�VhH�SpH�ChH�FpH�VpH�Cp�Fx�Sx�VxH���   �CxH���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   �SyH���   �Fy�Vy�Sz�Cy�Fz�VzH���   �CzH���   H����         H���   H���   H���   H���   ���   H���   ���   ���   ���   H��0[^_]A\Ð����H��(1�H�Q(H9Q sH����  �Phf���������H��(Ð���WVSH��0H�yHH��H�������������   H��H�\$(�C�������H�L$(�AX    Ɓ�    ����H�T$(1�H��f�ByH�BhH�B(    H�B     H�B0    H�BH�BH�B�B\�B`�Bd�b}��H��t@��H��uH��0[^_�1�H��0[^_�H��H��u�5� H���-}����� �#� �>� �[���H���1� H�L$(�W� H���/���H���鐐��������WVSH��@H��H��H����{ ���  H���{� H��H�KH���������   �{y ��   H���   H����  H��P(�����   �{y ��   H���   H����  H��P0����   H��twH�H���P0��u&�SXE1�A�   H�H�L$0�T$ H���P H�|$0�tDH���   H��@[^_À{z �h���H���   H��@[^_�fD  �{z t�H���r�������   1�H���   H��@[^_�f�     1�����f�     H���   H�SdH�CH+CH���   L�L���   H��I��H�D$ A�R8Hc�H�H���   H���   H)���   H���   H�C(    H�C     H�C0    H�H���   H�ChH���   H�CH�CH�C�C\�C`�Cd�����f�H�ChH�C(    H�C     H�C0    H�CH�CH�C����� H���   I���	'���l����7c �������WVSH�� H��H��L��H�IH�������uH��H	�uH�Cp   H��H�� [^_��     H��t�H��~�H��H�shH�{pH���       [^_Ð��ATUWVSH�� ���    H��H��L����   1�M��H�QH�A~	H9��k  H9�H���   ƃ�    ��H�Kh��D�cXH�PH���   H���   H�KH�CH�SH�{p�   HCCpH��H9�~$H���   H���`  H��P0A��t����   I��H��H�����  H�H��H�� [^_]A\Àyz u
D�aX1��f�H����  �Phf���t?H�Ch�Cz 1�D�cXH�C(    H�C     H�C0    H�CH�CH�C�M����     1��L�cH�SL9�t!I)�H��M��L��N%��L��LcH��H�H)�L�cH��     H�H)�t"H�<GI��H��L���Fy��H���taH��u�H��u&�Cy�����H��H���   f�W�H�P�x���H�ChH�C(    H�C     H�C0    �Cy H�CH�CH�C�����H� �Cb ��` ��������������UWVSH��8�AXH��H���   H��L��@��H���  H��P0����   @����   �{y uzL�C(H�C0L)�H���{z uH�SpH�J�H��HG�H=   �   HM�H9�BH�S H�t$ H�KHI��I)�I��L����y��H�H9�t<H��H)�H9Ÿ    HL�H��8[^_]ÐI��H��H��H��8[^_]��  f.�     �KXH�Sh��H�SH�SH�Su��t!H�KpH��vH�S(H�S H�TJ�H�S0�Cz�H�C(    H�C     H�C0    ���_ ���UWVSH��8H�����H��H��L���A    H��D���v�����uH��H��8[^_]�fD  H�NHA��H����w��H���t�1ҋ�$�   H�H��f�VyH���   H�F(    H�F     H�F0    H���   H���   H�Vh�~`�{H�      �VH�VH�VH��8[^_]Ð�����������AVAUATUWVSH��pH��H���   H��M��E��H����   H��    �P(��I�@��M��H�����L�sH���F    L��!�����<u@��tH��H��p[^_]A\A]A^�D  A��uzM��uu�{z tH���   H��P0��t^�C\1��{y �D$l��   �{z tH�{(H+{ H��1�A�   L���zv��H���t�HǋD$lH�>�F�{���f��   1��B���@ ���    t=H�C1�ƃ�    H9CH���   H�Kh��H�PH���   H���   H�KH�CH�SLcŋC\M�Ā{y �D$lu(�D$ H�L$PE��H�������H�D$PH��D$X�F�����A��uҋCdH�T$lH��L�D$8�D$l�/���L�D$8H�I��D$l멋CdH�T$lH�ىD$l����Hc���������UWVSH��HI�8I�hH�����H��H���A    H�JH�t�����tl���    t=H�C1�ƃ�    H9CH���   H�Kh��H�PH���   H���   H�KH�CH�SH�L$0�l$ E1�I��H�������H�D$0H��D$8�FH��H��H[^_]Ð�������VSH��X�AXH�ˉ���   �yy tw���    t=H�A1�H9AH���   ��H�PH���   H���   H�IhH�Cƃ�    H�SH�KH�SdH��������SdH�L$0A�   Lc��T$ H���6���H�|$0�t1H�S L�C(L9�s1f���tfA�0I��L�C(I)�H��I��������u]�����H��X[^ÐH�SpH����   f���f�t$Nu�Cz1�H��X[^�f.�     H�T$NA�   H���]�����t��Cz��멐�SXH�Ch��H�CH�CH�Cu��t#H�SpH��vH�C(H�C H�DP�H�C0�      �fD  H�C(    H�C     H�C0    f������i���H��X[^�D  �KXH�Ch��H�CH�CH�Ct8H�C(H�C H�DP�H�C0f����Cz�&���H�C(f�0H��H�C(��H��X[^Ð��u�H�C(    H�C     H�C0    뺐WVSH��@�AXH�ˉ��  �yz ��   H�AH;A���   ��   H�P�H�Q�P�1�f�����   f9����   @����   ���    H�Cu-H���   H�CH�S~H�Sƃ�   H���   H�C|H�CH�C�Cyf�0��H��@[^_�@ H����  �Phf���tsH�ChH�C(    ���   H�C     H�C0    �Cz H�CH�CH�CH�H�L$0H���D$    A�   I�������P H�|$0�tH�H���PHf��������������H��@[^_Ð��������������UWVSH��(�yX@��H��t~H�iHH��������tnH�^��H+^H���   H��H��t]H��P(��x��uH��H��([^_]��     H���r��H���   H��H��P@Hc�H��H�H��H�H��H��([^_]�H��������PX ����������������AUATUWVSH��X�AXH���  �yz �1  ���    H�A�j  H�SH9���  H���   �   H�{pHCspH��H�~���  H��P0���~  H���   H��P(����  Hc�H��H��H���   I��H���   H)�I)�H9�    LN��{y H���   tH�KH9K��  H9���  H��L���   ��  �C`M�L5 M��L���   L���   �Cd��  H�C1�M9�H�D$Hvr1�@ H���   L�D$HH�S`L�L�D$8L�xH�D$(H���   L�D$0M���      H�D$ A�R ������  H�D$HH+CI��I�����D  H����	����T  L���   A�   L��H+��   L�H;��   �T  H�KHM��L���~n��H����  H����s  1�H��   L���   I��H���   H�CM9�H�D$H�������Q  @���y���H�Ch��H�C(    H�C     H�C0    �Cy H�CH�CH�C��   H��� �\W H����  �Phf���t~H�ChH�C(    ���    H�C     H�C0    �Cz H�CH�CH�C�����1�H9Cƃ�    H���   H�Kh��H�PH���   H���   H�KH�CH9�H�S�a���� H��X[^_]A\A]�H�SH�KHI���@m��H��I����  H�ChH�C(    H�C     H�C0    �Cy H�CH�CH�C�����H��X[^_]A\A]�fD  L���   H�CH���   I)�L9�M��L��r0M��u1M��H���   �   ��	������f��   �=���fD  I��H��L�D- H���]��H���   H�붐H�� @���>���H�� ��U fD  M��~ZH�Ch�CXH�CH�Ct]J�`H�SH�C(    � H�C     H�C0    �Cy�����H���   H��P@H�H�l�H���R���@�������H�� �\U H�C�fD  H���X� H��I��u9H���   H��t�� L���   H���   �T���~��J���H��E1��� I��H���   I��L���U��� 1������H��t&H9��L���   E1�I��L���"��L���   �����H9�~�H����� I���i���H��� �T �(S ��������VSH��(H��H����  H�h� H�F@    H�H�CHH�      �FH�CP�FP�CXH�CH    �CP �CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �Fx�Cy�Cy �Fy�Cz�Cz �Fz�C|f�F|H���   Hǃ�       H���   H���   Hǃ�       H���   ���   ƃ�    ���   H���   H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H�ChH�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��([^Ð���������ATUWVSH�� L�%�8 I�D$H�q8H��H�H�A    H�{HH�A    H�A    H�A     H�A(    H�A0    H���a H�}� H��H�C@    H�H�S@�k��1�1��Cz H�CX    H��H�C`    H�Ch    H�Cp   f�Cxf�S|Hǃ�       Hǃ�       ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       �*g ��uH�� [^_]A\�H���w H���   H�� [^_]A\�H��H����j��I�T$H��H���` H����k����������������VSH��(H��H����  H�h� H�F@    H�H�CHH�FH�CP�FP�CXH�CH    �CP �CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �Fx�Cy�Cy �Fy�Cz�Cz �Fz�C|f�F|H���   Hǃ�       H���   H���   Hǃ�       H���   ���   ƃ�    ���   H���   H���   H���   Hǃ�       H���   H���   Hǃ�  �           H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H�ChH�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��([^Ð���������ATUWVSH�� L�%�5 I�D$H�q8H��H�H�A    H�{HH�A    H�A    H�A     H�A(    H�A0    H���^ H�}� H��H�C@    H�H�S@�h��1�1��Cz H�CX    H��H�C`    H�Ch    H�Cp   f�Cxf�S|Hǃ�       Hǃ�       ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       �*d ��uH�� [^_]A\�H���t H���   H�� [^_]A\�H��H����g��I�T$H��H���] H����h����������������SH�� H�t� H��H�����H�KH�g��H�4 H�K8H��H��] H��H�� [�<� ������������SH�� H�$� H��H��i���H�KH�Pg��H��3 H�K8H��H�H�� [�4] ����SH�� H�� H��H��)���H�KH�g��H��3 H�K8H��H�H�� [��\ ����VSH��(H��H�������H��H���D�  H�SHH�FHH�VH�SPH�CH�FP�VP�CP�CX�CX    �FX�C\�F\�C`�F`�Cd�FdH�ChH�Ch    H�FhH�CpH�Cp   H�Fp�Cx�Cx �FxH���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   H���   Hǃ�       H���   �Cy�Cy �Fy�Cz�Cz �FzH���   Hǃ�       H���   H���   Hǃ�       H���   ���   ƃ�    ���   H�Ch�      H�C(    H�C     H�C0    H�CH�CH�C�C\�C`�CdH��H��([^ÐSH�� H��H�I追��H��H�tHX�1�H��H�� [�& @ HX�S H�ك�H�� [�& ���������SH�� H�H��H�I�l���H��H�tHX�1�H��H�� [�a& �HX�S H�ك�H�� [�I& ���������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���#
 H���   H����" H���   H����" H���   H�OH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�U���   H�GH�WH�UH�EH��([^_]逽��SH�� H��H�I诿��H��t
H�� [�@ H�HX�S H�ك�H�� [�F% ������H��`������������ATUWVSH�� L�%'> H���   H��H��H��� 1�L�#H��f���  I�D$(H���   H�FHǃ�      Hǃ�      Hǃ�      H�CH�Hǃ�      Hǃ�      H�x�H�H���~ H���  H���! H���   H�VHǇ�       H���  ���   ���  ���   H�{Hǃ�      H�����  H�� H�F    H�H��PH���   H��(H�C�|���H���  H�� [^_]A\�H��H�01 H��H��H���   �- H���c��H�6= L�#H��H�KH�C    �Ð���������AVAUATUWVSH�� H�-�< H���   H��I��H��E���# 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    �c! L�%�< 1�H��I�D$(L��      cH���   �B! H�� H�H�{H��PH���   H��(H��H�C�����H��H���! E��L��H�������H�H�J�H�H��t!1��" �H�� [^_]A\A]A^�f.�     �Q ���" �H�� [^_]A\A]A^�I��H���
���L��L�cH�+H��H�C    H��/ H��H��H���   � H���b������H���Ր���������AVAUATUWVSH�� H�-#; H���   H��I��H��E��� 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    �� L�%�: 1�H��I�D$(L�cH���   � H�S� H�H�{H��PH���   H��(H��H�C�Y���H��H���~ I�U E��H���/���H�H�J�H�H��t 1��)! �H�� [^_]A\A]A^�f�     �Q ���! �H�� [^_]A\A]A^�I��H���z���L��L�cH�+H��H�C    H��- H��H��H���   �� H���s`������H���Ր���������AUATUWVSH��(H�-�9 H���   H��H��� 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    �K L�%l9 1�H��I�D$(L�cH���   �* H�ˡ H�H�{H��PH���   H��(H��H�C�����H��H���� �H��([^_]A\A]�H��H��, H��H��H���   �� H���S_��I��H������L��L�cH�+H��H�C    ����쐐�����������ATUWVSH�� H�BH��H��H�H�JH�P�L��H�I�PH�SH�h�I� H��      L�`�H��M�L���� H���   H���� I��$�   IǄ$�       H���   A��$�   ���   A��$�   Hǅ�       ���   H�F H�kH�G    H��H�CH�@�H�V(H�TH�FH�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�WH�C�����H�H�@�H���   H�� [^_]A\�H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    �]������ATUWVSH�� H�BH��H�H��H�JH�P�L��E��H�1�H�C    H�H�H��� H�F 1�H�CH�@�H�LH�F(H��� H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C�Q���H�H��H�H�H��o E��H��H���!���H�H�J�H�H��t1�� �H�� [^_]A\ËQ ��� �H�� [^_]A\�H��H���}���H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    �W\����ِ��ATUWVSH�� H�BH��H�H��H�JH�P�L��E��H�1�H�C    H�H�H�� H�F 1�H�CH�@�H�LH�F(H��b H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C�����H�H��H�H�H�� H�U E��H�������H�H�J�H�H��t1�� �H�� [^_]A\ËQ ��� �H�� [^_]A\�H��H������H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    ��Z����ِ��      UWVSH��(H�BH��H�H��H�JH�P�H�1�H�C    H�H�H��) H�F 1�H�CH�@�H�LH�F(H��
 H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C����H�H��H�H�H�� �H��([^_]�H�VH�H�R�H�NH�H��H�C    �Z��H��H�������H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�L��̐�������SH�� H�ܛ H�H��PH��H���   H�IH��(H�A�H��� H�����H�K`�_X��H��$ H�KPH��H�C�GN H�3 H�C    H�CH��2 H�H��& H���   H��H���   � H��H�� [鿑 ���������������SH�� H�,� H�H��PH��H���   H�IH��(H�A�H� � H��h���H�K`�W��H�$ H�KPH��H�C�M H�X2 H�C    H�CH��1 H�H�& H���   H��H���   H�� [� �������VSH��(H�H��H�H�@�H��H�R@H�IH�T�H�FHH�A�H�^� H��Ʋ��H�K`�W��H�v# H�KPH��H�C��L H�FH�H�@�H�V0H�H�F8H�CH�F H�CH�@�H�V(H�TH�FH�H�@�H�VH�H�C    H��([^Ð��UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H����� H���   H���� H���   H��� H���   H�MH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�W���   H�EH�UH�WH�G�h���H��H��([^_]Ð�����������SH�� H���      H�I����H��H�tHX�1�H��H�� [�4  @ HX�S H�ك�H�� [�  ���������SH�� H�H��H�I�<���H��H�tHX�1�H��H�� [�� �HX�S H�ك�H�� [�� ���������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���� H���   H��� H���   H��� H���   H�OH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�U���   H�GH�WH�UH�EH��([^_]�>�����������������SH�� H��H�I�_���H��t
H�� [�@ H�HX�S H�ك�H�� [� ������H��`�'����������ATUWVSH�� L�%/ H���   H��H��H���� 1�L�#H��f���  I�D$(H���   H�FHǃ�      ƃ�   Hǃ�      H�CH�Hǃ�      Hǃ�      Hǃ�      H�x�H�H����� H���  H��� H���   H�VHǇ�       H���  ���   f���  ���   H�{Hǃ�      H�����  H�ߖ H�F    H�H��PH���   H��(H�C�4���H���  H�� [^_]A\�H��H��! H��H��H���   �u H����S��H��. L�#H��H�KH�C    �Ð�AVAUATUWVSH�� H�-�- H���   H��I��H��E���s 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    �� L�%�- 1�H��I�D$(L�cH���   � H��� H�H�{H��PH���   H��      �(H��H�C����H��H���w E��L��H���y���H�H�J�H�H��t1��# �H�� [^_]A\A]A^� �Q ��� �H�� [^_]A\A]A^�I��H�������L��L�cH�+H��H�C    H�� H��H��H���   �� H���SR������H���Ր���������AVAUATUWVSH�� H�-, H���   H��I��H��E����  1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    �< L�%], 1�H��I�D$(L�cH���   � H�� H�H�{H��PH���   H��(H��H�C����H��H���� I�U E��H�������H�H�J�H�H��t1�� �H�� [^_]A\A]A^�f��Q ���u �H�� [^_]A\A]A^�I��H���Z���L��L�cH�+H��H�C    H�^ H��H��H���   �K  H����P������H���Ր���������AUATUWVSH��(H�-�* H���   H��H���[� 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    � L�%�* 1�H��I�D$(L�cH���   � H��� H�H�{H��PH���   H��(H��H�C����H��H���_ �H��([^_]A\A]�H��H�7 H��H��H���   �$� H���O��I��H�������L��L�cH�+H��H�C    ����쐐����ATUWVSH�� H�BH��H��H�H�JH�P�L��H�I�PH�SH�h�I� H�L�`�H��M�L���F� H���   H��� I��$�   IǄ$�  �           H���   A��$�   f���   A��$�   Hǅ�       ���   H�F H�kH�G    H��H�CH�@�H�V(H�TH�FH�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�WH�C����H�H�@�H���   H�� [^_]A\�H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    �N�����ATUWVSH�� H�BH��H�H��H�JH�P�L��E��H�1�H�C    H�H�H��Q H�F 1�H�CH�@�H�LH�F(H��2 H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C����H�H��H�H�H��� E��H��H�������H�H�J�H�H��t1�� �H�� [^_]A\ËQ ���t �H�� [^_]A\�H��H���]���H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    �L����ِ��ATUWVSH�� H�BH��H�H��H�JH�P�L��E��H�1�H�C    H�H�H��� H�F 1�H�CH�@�H�LH�F(H��� H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C����H�H��H�H�H�� H�U E��H������H�H�J�H�H��t1��* �H�� [^_]A\ËQ ��� �H�� [^_]A\�H��H�������H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�LH�VH�H�R�H�NH�H��H�C    �FK����ِ�UWVSH��(H�BH��H�H��H�JH�P�H�1�H�C    H�H�H�      �� H�F 1�H�CH�@�H�LH�F(H��z H�FH�{H��H�H�@�H�V0H�H�F8H�CH�H�H�@�H�V@H�H�FHH�C�Y���H�H��H�H�H��' �H��([^_]�H�VH�H�R�H�NH�H��H�C    �jJ��H��H������H��H�VH�H�R�H�N0H�H�V8H�SH�V H�SH�R�H�N(H�L��̐�������SH�� H��� H�H��PH��H���   H�IH��(H�A�H��� H������H�K`�H��H�( H�KPH��H�C�> H�x$ H�C    H�CH��# H�H�# H���   H��H���   �� H��H�� [�� ���������������SH�� H��� H�H��PH��H���   H�IH��(H�A�H�Њ H�����H�K`��G��H�x H�KPH��H�C��= H��# H�C    H�CH��" H�H�s H���   H��H���   H�� [�W� �������VSH��(H�H��H�H�@�H��H�R@H�IH�T�H�FHH�A�H�.� H��v���H�K`�]G��H�� H�KPH��H�C�E= H�FH�H�@�H�V0H�H�F8H�CH�F H�CH�@�H�V(H�TH�FH�H�@�H�VH�H�C    H��([^Ð��UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���C� H���   H���d H���   H���U H���   H�MH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�W���   H�EH�UH�WH�G�F���H��H��([^_]Ð���������VSH��   E1�H��H��H�L${H���1$  �|${ t~H��D$|    H�P�H��      H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R`�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �� H��H�Ĉ   [^��* H��H��t �=� H�H�p�HރN �Fu7�D� ��� H�HX�K �Cu跇 貇 H���� H���"F��蝇 H���� H���F���������������VSH��   E1�H��H��H�L${H����"  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R�T$|��uH��H�Ĉ   [^�H�H�H�H�Q � H��H�Ĉ   [^��[) H��H��t �� H�H�p�HރN �Fu7�� ��� H�HX�K �Cu�g� �b� H���ʁ H����D���M� H��赁 H���D���������������VSH��   E1�H��H��H�L${H���!  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�RP�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �M H��H�Ĉ   [^��( H��H��t �~ H�H�p�HރN �Fu7褀 ��}~ H�HX�K �Cu�� �� H���z� H���C����� H���e� H���mC���������������VSH��   E1�H��H��H�L${H���A   �|${ t~H��D$|    H�P�H�H��H�� �        H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�RX�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �� H��H�Ĉ   [^��& H��H��t �M} H�H�p�HރN �Fu7�T ��-} H�HX�K �Cu�ǃ � H���* H���2B��譃 H��� H���B���������������VSH��   E1�H��H��H�L${H����  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�RH�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �
 H��H�Ĉ   [^��k% H��H��t ��{ H�H�p�HރN �Fu7�~ ���{ H�HX�K �Cu�w� �r� H����} H����@���]� H����} H����@���������������VSH��   E1�H��H��H�L${H���  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R(�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �]	 H��H�Ĉ   [^��$ H��H��t �z H�H�p�HރN �Fu7�| ��z H�HX�K �Cu�'� �"� H���| H���?���� H���u| H���}?���������������VSH��   E1�H��H��H�L${H���Q  �|${ t~H��D$|    H�P�H�H��H��   H�����         L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R�T$|��uH��H�Ĉ   [^�H�H�H�H�Q � H��H�Ĉ   [^���" H��H��t �]y H�H�p�HރN �Fu7�d{ ��=y H�HX�K �Cu�� �� H���:{ H���B>��� H���%{ H���->���������������VSH��   E1�H��H��H�L${H���  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R0�T$|��uH��H�Ĉ   [^�H�H�H�H�Q � H��H�Ĉ   [^��{! H��H��t �x H�H�p�HރN �Fu7�z ���w H�HX�K �Cu�~ �~ H����y H����<���m~ H����y H����<���������������VSH��   E1�H��H��H�L${H���  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R �T$|��uH��H�Ĉ   [^�H�H�H�H�Q �m H��H�Ĉ   [^��+  H��H��t �v H�H�p�HރN �Fu7��x ��v H�HX�K �Cu�7} �2} H���x H���;���} H���x H���;���������������VSH��   E1�H��H��H�L${H���a  �|${ t~H��D$|    H�P�H�H��H��   H����   L��� �        H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R8�T$|��uH��H�Ĉ   [^�H�H�H�H�Q � H��H�Ĉ   [^��� H��H��t �mu H�H�p�HރN �Fu7�tw ��Mu H�HX�K �Cu��{ ��{ H���Jw H���R:����{ H���5w H���=:���������������VSH��   E1�H��H��H�L${H���  �|${ t~H��D$|    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�t$0H�D$@    H�D$H��  L�D$PL�D$|L�D$(L�D$PH�D$ A�R@�T$|��uH��H�Ĉ   [^�H�H�H�H�Q �� H��H�Ĉ   [^�� H��H��t �t H�H�p�HރN �Fu7�$v ���s H�HX�K �Cu�z �z H����u H���9���}z H����u H����8���������������WVSH�� H�H�@�H��H��L��H���   H��t$H��
   �PPI��H��H��D��H�� [^_�   �� ���ATUWVSH��0H��H�A    H��L��H�L$/A�   H��E���_  �|$/ u(H�NH��~E1�fD�H���O  H��H��0[^_]A\ÐH�H�@�H���   H�CH9Cwr�    H�H���PHH�NH�QH9�|ef.�     f���u�H��~f�  H�ɺ   ��   �   ��   �     �H��H�Sf���tSH�CH;Cs�H�N� H�QH9�}�f�����   fD9���   H��f�G�H�VH�SH;Sr�H�H���PPf���u�H��H�F��   1�H��f��   uU���PH���      H����   ��q H�H�H�H�I �A��   ��s H����   H�~ f�  ����� �   H�H�H�H�Q �9  H��H��0[^_]A\�1�H��~f�  H���v�����u�H��H��0[^_]A\�@ H��������   ��뢺   ��Qq H�Hp�N �Ft��w ��w H���Ns H���V6����w H�N� ���H���0s H���86����������VSH��(H�H�@�H��H��H���   H��t H��
   �PPH��H��D��H��([^�   � �����������ATUWVSH��0H��H�A    H��E��H�L$/D��H��A�   �  �|$/ ��   H�H�@�H���   H�CH9C��   � f�����   fD9�uK�ef�f�H��H�O(H�FH�SH;S��   �H��H�Sf���taH�CH;Csw� f���tNf9�tH�O(H;O0r���H�H���Phf���u�H�~ u�   H�H�H�H�Q �O� H��H��0[^_]A\ÐH�~҃����АH�H���PP�{���f�H�H���PH�~���f�H�H���PH����H��H��u�do H�Hp�N �Ft#��u �Io H�H�x�H��O �Gt��u ��u H���Cq H���K4���6q H�~ �5����G���H���q H���&4��������VSH��8A�   H��H�A    H��H�L$/H����  �|$/ u2H�{ u�   H�H�H�H�Q �4� H��H��8[^�f.�     H�H�@�H���   H�QH9Qv7�H��H�Qf���tH�C   f�H��H��8[^ÐH�{҃���닐H��PP��H��H��u�*n H�HX�K �Ct#��t �n�       H�H�p�HރN �Ft�t �t H���	p H���3����o H�{ �����(���H����o H����2��������������SH��0A�   H��H�A    H�L$/H���  �|$/ ��   H�H�@�H���   H�QH9Q��   �H��H�Qf���tH�C   H��0[�fD  H�{҃���H�HX�S H���� �����H��0[�H��H��t8�m H�H�P�HڃJ �BuO�o H�{ uǺ   뮐H��PP�{�����l H�HX�K �Ct�js �es H����n H����1���Ps H���n H����1������������������SH��@A�   H��H�A    H�L$?H���  �|$? tLH�H�@�H���   H�AH9Av]� f���t5H��@[�H��H��tM� l H�HX�K �Cug�*n �����H��@[�H��D$,HZ�S H�ك��v� �D$,�H��PH���k H�HX�K �Ct�mr �hr H����m H����0���Sr H���m H����0�����WVSH��0H��H�A    H��L��H�L$/A�   H���  �|$/ t$H�I��H��H�@�H���   H��P@H9�H�CuH��H��0[^_�H�H�H�HًQ ���� H��H��0[^_�H��H��t �k H�H�x�H߃O �Gu7�m ���j H�HX�K �Cu�{q �vq H����l H����/���aq H����l H����/���UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H����� H���   H���� H���   H���� H���   H���   H���   ���   H���   ���   f���   ���   f��� �        ���   ���   H�W���   H�EH�UH�GH��([^_]Ð���������SH��@A�   H��H�L$?H����  �|$? tNH�H�@�H���   H��t:H��P0���t61�H��@[�H��H��tD�i H�HX�K �Cu^�k  �������H��D$,HZ�S H�ك���� �D$,��Ei H�HX�K �Cu��o ��o H���Bk H���J.����o H���-k H���5.�������SH��`)|$PH��o:H��H�H�HًQ ����j� H�L$OA�   H����
  �|$O t:H�H�P�H��B u*H���   H�L$0)|$ A�   L�D$ H��P(H�|$0�t(|$PH��H��`[��     H�H�H�HًQ ����� ��H��H��t �Kh H�H�H�HكI �Au7�Rj ��+h H�HX�K �Cu��n ��n H���(j H���0-���n H���j H���-�������������WVSH��PH�H��H�H�H��D��HًQ ����K� H�L$OA�   H����	  �|$O t8H�H�P�H��B u(H���   H�L$0A��I��H��D$    �P H�|$0�tH��H��P[^_�H�H�H�HًQ ����� ��H��H��t �9g H�H�p�HރN �Fu7�@i ��g H�HX�K �Cu�m �m H���i H���,���m H���i H���	,�����������VSH��XA�   H�����H��H���A    H�L$O��  �|$O tBH�H�P�H��B u2H���   H�L$0A�   E1�H��D$    �P H�D$0H��D$8�CH��H��X[^�H��H��t�Ef H�Hp�N �Fu7�Oh ���(f H�Hp��      N �Fu��l �l H���%h H���-+���l H���h H���+����������SH��0H�H��H�A    H�H�HًQ ����K� H�L$/A�   H����  �|$/ t2H�H�H�H�H���   H��t5H�PH9PsAH�J�H�H�B�f���tH��H��0[�fD  H�H�H�HًQ ����� H��H��0[�f�L� ���  H��A�PX�H��H��u�!e H�HX�K �Ct#�k �e H�H�P�HڃJ �Bt�k �k H��� g H���*����f �_���H����f H����)����������������SH��0A�   H��H�A    H�L$/H���  �|$/ t2H�H�@�H���   H�QH9Qv"�H��H�Qf���tH�C   H��H��0[�H��PP�� H�H�H�HًQ ���� H��H��0[�H��H��u�d H�HX�K �Ct#�j ��c H�H�P�HڃJ �Bt�j �j H����e H����(����e �m���H����e H����(���AVAUATUWVSH��0H��H��H���4  H�A    A�   H��H�L$/�  H����   �l$/@����   H�H�@�H���   H�GH9G�t  � H�SE1�I��������I�       �D  H9�~Rf�����   L�OI��H�OI)�L��H)�H��L9�IO�H����   H�AH�I9�H�OH�S��   H9���L9���   f���tL�kA��H�       ���    E��tH��������H�CH�H�H�HًQ ���� �     H��H��0[^_]A\A]A^�����H��0[^_]A\A]A^�f.�     H��������H9�t�E��t�H�C�      �fD  H��I9�H�Sv9�H��H�Of���t�H�GH;Gs� H�S�����H�H���PHH�S����H�H���PP��H�H���PH����E��tL�sf���>�������H��H��u�a H�HX�K �Ct#�5h �a H�H�x�H߃O �Gt�h �h H���zc H���&���mc H�������H���]c H���e&�������AWAVAUATUWVSH��8fA���H��H��D��D���}  H�A    A�   H��H�L$/�  H���E  D�l$/E���6  H�H�@�L���   I�D$I9D$�*  � H�KE1�I�       � H9�~f����  f9���   M�T$I��M�L$I)�L��L)�H��L9�LN�I���!  M��M��tL��L��f98��   H��H��u�K�YL�I9�I�D$H�K��  H9�� �H��������H9��  f�����   f9���  L�{E��H�       ��@���H��������H9��m  E����   H��H�KI�D$I;D$�=  H��I�D$ H��H��8[^_]A\A]A^A_��������D  H��������H9�tqE��tH�CH�H�H�HًQ ����� H���L)�H��I��I��� ���H��M9�H�K��   A�I��M�L$f���t�I�D$I;D$sm� H�K�a����E��t�H��������H�C�E��tfD  H��������H�{f����`���f9�����H�KH��������H9����������� I�$L���PHH�K�����I�$L���PH�����I�$L���PP�P���I�$L���PP�����E���w����E��t��k���H��H��u�=^ H�HX�K �C�      t#��d �"^ H�H�x�H߃O �Gt�d �d H���` H���$#���` H���J���H����_ H���#���������UWVSH��(H�H��� H�H�H��D��HыQ ����   H���   H����   H����  H�H�H�H���  �A�  H���   H�CH;C�  � H���   H���#  f���u-�m �H��H�Sf���tOH�CH;C��   � f���t8L�M D���    H��A�Q����   H�SH;Sr�H�H���PPf���u� H�Hp�H��Q ����H��([^_]�P� E��u
�A�>����H��([^_]�H��H��ty�\ H�H�X�H�K �C��   �^ f.�     H�Hp�H��Q ��t���H��([^_]��� H�H���PH�#����H�H���PHH�H�J�H������� �\ H�Hp�N �Ft�b �b H���^ H���#!���b H���^ H���!����������������UWVSH��(H�H��� H�H�H��D��HыQ ����   H���   H����   H����  H�H�H�H���  �A�  H���   H�CH;C�  � H���   H���#  f���u-�m �H��H�Sf���tOH�CH;C��   � f���t8L�M D���    H��A�Q����   H�SH;Sr�H�H���PPf���u� H�Hp�H��Q ����H��([^_]�P� E��u
�A�>����H��([^_]�H��H��ty�Z H�H�X�H�K �C��   �\ f.�     H�Hp�H��Q ��t���H��([^_]��� H�H���PH�#����H�H���P�      HH�H�J�H������� �Z H�Hp�N �Ft�` �` H���\ H���#���` H���\ H�������������������WVSH�� H�H�@�H��H��L��H���   H��t$H��
   �PPI��H��H��D��H�� [^_�   �� ���AWAVAUATUWVSH��8H��H�A    H��M��H�L$/A�   H��E��D���v����|$/ �  H�H�@�H���   H�FH9F��  � L�OI�IL9���   f�����  f9�L�VH�V�  M��M)�M�F�M��I)�I��M9�MN�I���;  H��M��tH��L��f9�	  H��H��u�O�< H��M�������L�OL�VH�VL�M�L�L9�H�VL�O�%  I�I�L9��[���f�����  fD9��l  M���G  1ɺ   f�M �$H�H���PPf�M��H�O~c1�H��f�U u]�   H�H�H�H�Q �� �DI��H��H���k  ��W H�H�p�H��N �F�i  ��Y M���`  H�OH��t�H��H��8[^_]A\A]A^A_�H)�I��I��I��M������������f�E L�uI9�H�Ovs�H��H�Vf���t:H�FH;Fsj� L��L�O�>���D  H�H���PH�'���H�H���PH����L�OL��M��   ~1�f�E M��������������H�H���PP덺   ��H�H���PHL�OL�������L�VH�VI9�H�O�����H��M��H�V����������M��~E1�I���fD�E ���������   �u������������V H�Hx�O �Gt5�] �] H� fA�  �;�������H���jX H���r���:�      �����\ H���PX H���X����������VSH��8H�H��H�A    H�H��HًQ ����� H�L$/A�   H�������|$/ t7H�H�H�H�L���   M��t5I�HI9Hs@�A�f9�u7H��I�Hf���t
H��H��8[^�H�H�H�HًQ ���� H��H��8[^�I� ��L���PX��H��H��u�bU H�HX�K �Ct#��[ �GU H�H�p�HރN �Ft��[ ��[ H���AW H���I���4W �h���H���'W H���/�����������������WVSH��0H��H�A    H��L��H�L$/A�   H��������|$/ ��   H�H�@�H���   H�AH�QH9���   H)�H��H��~bH�H9�HN�I��H�R�H���   H��L�	A�Q@H�CH��0[^_�H��H��tR�RT H�H�x�H߃O �Gui�YV H�CH��0[^_�H���u�H�H�H�HًQ ���� ��H��P8�q���� T H�HX�K �Ct�Z �Z H����U H������Z H����U H����������������������UWVSH��(H�iH��H��H���� 1�H��Hǃ�       f���   H��[ H�H��(H�CH�Gƃ�    Hǃ�       Hǃ       H�CH�Hǃ      Hǃ      H�p�H�H���p� H���   H����� H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   H�G    H��([^_]�H��H�g� H��H�PH�S�W� H���������������������WVSH�� H�qH��H��H���w� 1�H��H��f���   H��Z H�H��(Hǃ�       ƃ�    �      Hǃ�       Hǃ       Hǃ      Hǃ      H�CH�C    ��� �H�� [^_�H��H��� H��H�PH�S�� H���������������������WVSH�� H�qH��H���� 1�ƃ�    1�f���   H��H��Y Hǃ�       H�H��(Hǃ�       Hǃ       Hǃ      Hǃ      H�CH�C    �� �H�� [^_�H��H��� H��H�PH�S��� H���T������WVSH�� H�L��H�L�BH�P�L�H�WH�QHH�H�H��H�p�H�H���3� H���   H���� H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   H�G    H�� [^_Ð����H�H�L�JH�P�L�L��H�A    HH��� ����������H�H�L�BH�P�L�1�H�A    HH���� �����������SH�� H�\X H�H��� H��H�A    H�IH��H��� H��H�� [�M ��H�!X H�H�� H��H�A�    H��H��g� �������H�H�H�@�H�RH�H�A    Ð����UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���� H���   H���� H���   H����� H���   H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�U���   H�GH�WH�EH��H��([^_]Ð������H�␐�����������SH�� H�H��H�H�H���H��H�� [Ð��SH�� H�H��H�H�H���H��H�� [Ð��VSH��8E1�H��H��H�L$.H�������|$. tBH�H�H�H�H���      tBH���   L�D$/H����� H���T$/t@��tH��   H�H�H��H��t=H��H��8[^ú   Q �� H��H��8[^�D  H�H�H�Hـ�҃������H��   H�H�H���H��H��t �M H�H�p�HރN �Fu7��O ��M H�HX�K �Cu�4T �/T H���O H������T H���O H����������������+���������������k����������������������������������������������+��������������VSH��   E1�H��H��H�L$wH�������|$w ��   H��D$x    H�P�H�H��H��   H����   L���   H�L$`H�D$X��  L�L�L$@H�D$ H�D$@    H�D$H��  L�D$PL�D$|L�D$0L�D$xL�D$(L�D$PA�R�D$|��T$x��uH��H�Ĉ   [^�H�H�H�H�Q �� H��H�Ĉ   [^��|� H��H��t �L H�H�p�HރN �Fu7�N ���K H�HX�K �Cu�R �R H����M H�������nR H����M H������������������������������������K�����������������������������VSH��   E1�H��H��H�L$wH�������|$w ��   H��D$x    H�H�H�H��   H��H����   L���   L�L$@H�D$X��  L�H�L$`H�D$@    H�D$H��  H�D$ L�D$PL�D$|L�D$0L�D$xL�D$(L�D$PA�R�D$|�T$x= ���} ��� ����T$xf���u'H��H�Ĉ   [^�=�  ~5����  �҉T$xf�t�H�H�H�H�Q � � H��H�Ĉ   [^� f�����       H��H��t'�HJ H�H�p�HރN �Fu>�OL �T$x�y����!J H�HX�K �Cu�P �P H���L H���&���P H���	L H�������;���������������{�����������������������������UWVSH��8H�|$ H�ΉӉ�H��H���  �|$  t*H�H�@�H���   H�A(H;A0sqf�H��H�A(f���tAH�D$(H�HB��@ H��t ��� ��uH���   H��tH��P0���t;H��H��8[^_]�H�H�H�H�Q ���� ��     H����Ph��� H�L$(H�HH�Q ���i� �H��H��u.��H H�Hp�N �Ft6�cO H��H���  H�������H H�H�X�H�K �Ct�2O �-O H���J ���J �	���H���J 믐��������������VSH��(H�HH�H�H��H�X�H�H��讱 H���   H����� H���   H����� H���   H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   ���   H��([^Ð������SH�� H�H�@�H��H���   H��tH��P0���t	H��H�� [�H�H�H�HًQ ����� H��H�� [�H��H��t �TG H�H�P�HڃJ �Bu7�[I ��4G H�HX�K �Cu��M ��M H���1I H���9���M H���I H���$������SH��@H�L�
L�RH��H�H�H��A u/H���   L�D$ L�L$ A�   H�L$0L�T$(H��P(H�|$0�tH��H��@[�f�     H�H�H�HًQ ���� H��H��@[�H��H��t �dF H�H�      �P�HڃJ �Bu7�kH ��DF H�HX�K �Cu��L ��L H���AH H���I����L H���,H H���4������SH��@H�H��H�H�H��A u,H���   H�L$0E��I��L�H���D$    A�R H�|$0�tH��H��@[� H�H�H�HًQ ���+� H��H��@[�H��H��t �E H�H�P�HڃJ �Bu7�G ��dE H�HX�K �Cu��K ��K H���aG H���i
����K H���LG H���T
������VSH��HH�H��H�����H���A    H�H�H��A u2H���   A�   E1�H�L$0H��D$    �P H�D$0H��D$8�CH��H��H[^�H��H��t�D H�Hp�N �Fu7�F ���D H�Hp�N �Fu�)K �$K H���F H���	���K H���wF H���	�����������������UWVSH��8H�\$ H��H��H��H��L���/  �|$  t H�I��H��H�@�H���   H��P`H9�uHH�D$(H�HB��@ H��t �� ��uH���   H��tH��P0���t3H��H��8[^_]��    H�H�H�H�Q ���+� �f�     H�L$(H�HH�Q ���	� �H��H��u�iC H�Hp�N �Ft#�J �NC H�H�x�H��O �Gt"��I ��I H���HE H���  H���H���3E ����H����H���!E �א��������������SH��0H�H��� H�QH�H�H�H��H���   D�@ H��t5E��tD��H����H��0[�<� H�T$(�����H�T$(H�HP�D�B H��E��u��H��0[ÐSH��0H�H��� H�QH�H�H�      �H��H���   D�@ H��t5E��tD��H����H��0[��� H�T$(����H�T$(H�HP�D�B H��E��u��H��0[ÐVSH��(H�AH�H��HB��@ H��t �� ��uH���   H��tH��P0���tH��([^�H�NH�HH�Q ��H��([^�@� VSH��(H�AH�H��HB��@ H��t �>� ��uH���   H��tH��P0���tH��([^�H�NH�HH�Q ��H��([^��� VSH��(H�H�@�H��L��H���   H��P`H9�u
H��([^� H�HX�S H�ك�H��([^�� �����ATUWVSH��`H�l$PH��I��H��H��������|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@L�d$(�D$ M��L�D$0L�D$0��H�T$8H��A�RH�|$H tH�H�H�H�Q ����� H�D$XH�HB��@ H��t ��� ��uH���   H��tH��P0���tKH��H��`[^_]A\�f�     H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��%���H�L$XH�HH�Q ���E� ��� �	� H��H��u.�? H�Hp�N �Ft6�5F H��H���j���H������m? H�H�x�H��O �Gt�F ��E H���gA ���`A �����H���SA 믐ATUWVSH��`H�l$PH��A��H��H��� ����|$P ��   H�H�X�H�H���   H���  ���    E����   ���   L�A�    ��H��L���   H�L$@D�d$(�D$ M��L�L$0I��A��L�D$8L�D$0A�R�|$H tH�H�H�H�Q ���� H�D$XH�      �HB��@ H��t �� ��uH���   H��tH��P0���tEH��H��`[^_]A\� H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��)���H�L$XH�HH�Q ���u� ��>� �9� H��H��u.��= H�Hp�N �Ft6�eD H��H������H�������= H�H�x�H��O �Gt�4D �/D H���? ���? �����H���? 믐UWVSH��x)t$`H�l$PH��H��H��f(��L����|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@�D$ �t$(M��L�D$0L�D$0��H�T$8H��A�R8�|$H tH�H�H�H�Q ���7� H�D$XH�HB��@ H��t �=� ��uH���   H��tH��P0���tF(t$`H��H��x[^_]ÐH���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��)���H�L$XH�HH�Q ���� ��n� �i� H��H��u.��; H�Hp�N �Ft6�B H��H�������H�������; H�H�x�H��O �Gt�dB �_B H����= ����= �����H���= 믐UWVSH��   �*�|$0H�l$pH��H��H���|����|$p ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$`�D$ �l$0M��L�D$P�|$@L�D$P��H�T$XH�T$@H�T$(H��A�R@�|$h tH�H�H�H�Q ���[� H�D$xH�HB��@ H��t �a� ��uH���   H��tH��P0���tJH��H�Ĉ   [^_]��    H���   H�      ��tFH��    �PPH�f���   ƃ�   H�Z�H�����H�L$xH�HH�Q ����� ��� �� H��H��u.�: H�Hp�N �Ft6�@ H��H�������H���"�����9 H�H�x�H��O �Gt�@ �@ H����; ����; �����H����; 믐ATUWVSH��`H�l$PH��A��H��H�������|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@D�d$(�D$ M��L�D$0L�D$0��H�T$8H��A�R�|$H tH�H�H�H�Q ���� H�D$XH�HB��@ H��t �� ��uH���   H��tH��P0���tKH��H��`[^_]A\�f�     H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��%���H�L$XH�HH�Q ����� ��� �� H��H��u.�K8 H�Hp�N �Ft6��> H��H������H���R����8 H�H�x�H��O �Gt�> �> H���: ���: �����H���: 믐ATUWVSH��`H�l$PH��A��H��H��������|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@D�d$(�D$ M��L�D$0L�D$0��H�T$8H��A�R �|$H tH�H�H�H�Q ���� H�D$XH�HB��@ H��t ��� ��uH���   H��tH��P0���tKH��H��`[^_]A\�f�     H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��%���H�L$XH�HH�Q ���%� ���� ��� H��H��u.�      �{6 H�Hp�N �Ft6�= H��H���J���H�������M6 H�H�x�H��O �Gt��< ��< H���G8 ���@8 �����H���38 믐ATUWVSH��`H�l$PH��I��H��H��� ����|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@L�d$(�D$ M��L�D$0L�D$0��H�T$8H��A�R(�|$H tH�H�H�H�Q ����� H�D$XH�HB��@ H��t ��� ��uH���   H��tH��P0���tKH��H��`[^_]A\�f�     H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��%���H�L$XH�HH�Q ���U� ��� �� H��H��u.�4 H�Hp�N �Ft6�E; H��H���z���H�������}4 H�H�x�H��O �Gt�; �; H���w6 ���p6 �����H���c6 믐ATUWVSH��`H�l$PH��I��H��H���0����|$P ��   H�H�X�H�H���   H���  ���    ��   ���   L��    ��I��L���   H�L$@L�d$(�D$ M��L�D$0L�D$0��H�T$8H��A�R0�|$H tH�H�H�H�Q ���� H�D$XH�HB��@ H��t �"� ��uH���   H��tH��P0���tKH��H��`[^_]A\�f�     H���   H��tFH��    �PPH�f���   ƃ�   H�Z�H��%���H�L$XH�HH�Q ���� ��N� �I� H��H��u.��2 H�Hp�N �Ft6�u9 H��H������H��������2 H�H�x�H��O �Gt�D9 �?9 H���4�       ���4 �����H���4 믐WVSH�� H�yH��H��H���W� 1�H��Hǃ�       f���   H��: H�H��(H�CH�ƃ�    Hǃ�       Hǃ�       Hǃ       Hp�Hǃ      H���<� H���   H��荽 H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   H�� [^_�H��H�<� H��H�PH�S�,� H����������WVSH�� H�qH��H��H���W� 1�H��H��f���   H��9 H�H��(Hǃ�       ƃ�    Hǃ�       Hǃ�       Hǃ       Hǃ      H�C賽 �H�� [^_�H��H��� H��H�PH�S耥 H���������������SH�� H��H�I诤 1�ƃ�    f���   H�09 H�H��(Hǃ�       Hǃ�       Hǃ�       Hǃ       Hǃ      H�CH�� [�WVSH�� H�qH��H���:� 1�ƃ�    1�f���   H��H��8 Hǃ�       H�H��(Hǃ�       Hǃ�       Hǃ       Hǃ      H�C藼 �H�� [^_�H��H�t� H��H�PH�S�d� H�������������������VSH��(H�H�HH�H�BH��H�I� H�p�L�H���ė H���   H���� H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   H��([^Ð��������������L�
L�	II�H�BL��H�鷻 �������H�H�H�@�H�RH�Ð������������H�H�HH�H�B1�H��x� ��������SH�� H�<7 H�H�J� H��H�IH���      H��7� H��H�� [�:, ����������H�7 H�H�� H��H��H���� ���������������H�H�H�@�H�RH�Ð������������WVSH�� H�H�p�H��H�H�H�X�H��H�H���w� H���   H��蘹 H���   H��艹 H���   H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   ���   H��H�� [^_Ð�����������H�␐�����������SH�� H�H��H�H�H���H��H�� [Ð��SH�� H�H��H�H�H���H��H�� [Ð�����������������WVSH��@H�|$0H��H��H��H�������|$0 t<H�H�H�H�H��trH���   L�D$/H���� H��uH��   H�H�H��M H��thH�D$8H�HB��@ H��t �A� ��uH���   H��tH��P0���tH��H��@[^_ú   Q �� �H�L$8H�HH�Q ���պ ��H��   H�H�H���H��H������H���O���H��H��u�, H�Hp�N �Ft-�2 ��+ H�H�X�H�K �Ct�2 ��- �(����~2 H����- �H����- 닐������������x������������;��������������H��8�*�|$ H�T$ �����H��8Ð�������Z����������������������������k������������������������������K��������������H�H�@�D��J��@t��t���P������H��������������������������������������������������������VSH��8H��H��H��n H����4���q  ��uA���         � �L������1�i�e�lЉ�H��H��p  u�Hǃ�	  p  H��8[^�H�6H�T$(E1�H��������> ��t
H�D$(�8 t�H��m �[� �����������WVSH�� H��H��H��m H���44����u4���Genuu��ubH�=mm H��m H��蔗��H��H�t1H�� [^_�H�Gm H��H�;��3����t�H�Fm H����3����t�H�Dm ��� �    H�=m �   ���   @t�H�    띐VSH��8H��� H��H�L�D$/H��H�I�����H��8[^�H��H��訽 H���`�������������������VSH��(H�C� H��H�L�BH��H�H�I�9����H��([^�H��H���V� H��������������������H��� H��H�H��H������������VSH��(H��1 H��H�H�I�Բ���H��([^�H��H���� H���������������SH�� H���   H��H�� [�& ������SH��0H�$1 H�H��H�I�������A���~H��蔼 �H��0[�H�T$/H�������H���w� �H��0[�SH�� H��H��H�I軥��H��H�� [Ð�SH�� H��A��H�I�+D��H��H�tHX�1�H��H�� [� � HX�S H�ك�H�� [�	� ���������SH�� H�H��A��H�I��C��H��H�tHX�1�H��H�� [�ͬ HX�S H�ك�H�� [鶬 ������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H��蓐 H���   H���d� H���   H���U� H���   H�OH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�U����         H�GH�WH�UH�EH��([^_]��C��SH�� H��H�I�F��H��t
H�� [�@ H�HX�S H�ك�H�� [鶫 ������H��X�GN���������ATUWVSH�� L�%W� H���   H��H��H���
� 1�L�#H��f���  I�D$(H���   H�FHǃ�      Hǃ�      Hǃ�      H�CH�Hǃ�      Hǃ�      H�x�H�H���� H���  H���� H���   H�VHǇ�       H���  ���   ���  ���   H�{Hǃ�      H�����  H�W. H�F    H�H��(H���   ��W��H���  H�� [^_]A\�H��H��� H��H��H���   襙 H������L�#H��H�C    �ΐ������������AUATUWVSH��(H�-�� H���   H��I��H��E��襘 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    �� H�V- H�H�{H��(H���   H���X��H��H��蹧 E��L��H��A���g@��H�H�J�H�H��t1��a� �H��([^_]A\A]� �Q ���E� �H��([^_]A\A]�I��H���\��L��H�+H��H�C    H�D� H��H��H���   �A� H��������H���א�AUATUWVSH��(H�-�� H���   H��I��H��E���U� 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    蕦 H�, H�H�{H��(H���   H���DW��H��H���i� I�$E��H��A���?��H�H�J�H�H��t�      1��� �H��([^_]A\A]�f��Q ����� �H��([^_]A\A]�I��H���l[��L��H�+H��H�C    H��� H��H��H���   �� H���i�����H���א�ATUWVSH�� H�-W� H���   H��H���� 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   H�C    �M� H��* H�H�{H��(H���   H����U��H��H���!� �H�� [^_]A\�H��H�� H��H��H���   �� H������I��H���EZ��L��H�+H��H�C    ����ATUWVSH�� H�BH��H�I��H�JH�P�L��H�I�PH�SH�x�I� H�H�h�H��L�H���6� H���   H���7� H���   Hǅ�       H���   ���   ���   ���   HǇ�       ���   I�$H�{H�F    H��H�H�@�I�T$H�H�V�=S��H�H�@�H���   H�� [^_]A\�I�T$H�H�R�I�L$H�H��H�C    �^�����������������ATUWVSH�� H�BH��H�H��H�JH�P�H�{L��E��H�1�H�C    H�H�H��}� H�H��H�H�@�H�VH��3T��H�H��H�H�H��Q� E��H��H��A����;��H�H�J�H�H��t1���� �H�� [^_]A\ËQ ���� �H�� [^_]A\�H��H���[X��H��H�VH�H�R�H�NH�H��H�C    �e����ې��ATUWVSH�� H�BH��H�H��H�JH�P�H�{L��E��H�1�H�C    H�H�H�荢 H�H��H�H�@�H�VH��CS��H�H��H�H�H��a� H�U E��H��A���;�      ��H�H�J�H�H��t1��� �H�� [^_]A\ËQ ���� �H�� [^_]A\�H��H���jW��H��H�VH�H�R�H�NH�H��H�C    �t����ې�UWVSH��(H�BH��H�H��H�JH�P�H�{H�1�H�C    H�H�H�襡 H�H��H�H�@�H�VH��[R��H�H��H�H�H��y� �H��([^_]�H�VH�H�R�H�NH�H��H�C    �����H��H���V��H���͐�����������SH�� H��& H�H��(H��H���   H��# H�AH�I�=��H�KX�V���H��� H�KHH��H�C�>�  H�o� H�C    H�H�ů H���   H��H���   辑 H��H�� [�� �SH�� H�& H�H��(H��H���   H�# H�AH�I�<��H�KX�����H�/� H�KHH��H�C��  H�߼ H�C    H�H�5� H���   H��H���   H�� [�)� ���������VSH��(H�H��H�H�@�H��H�RH�IH�T�H��" H���;��H�KX�5���H��� H�KHH��H�C��  H�FH�H�@�H�VH�H�C    H��([^Ð����������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���C� H���   H���� H���   H���� H���   H�MH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�W���   H�EH�UH�WH�G�T��H��H��([^_]Ð�����������SH�� H��A��H�I��Z��H��H�tHX�1�H��H�� [逩 HX�S H�ك�H�� [�i� ���������SH�� H�H��A��H�I�Z���      H��H�tHX�1�H��H�� [�-� HX�S H�ك�H�� [�� ������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���Ӄ H���   H����� H���   H���� H���   H�OH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�U���   H�GH�WH�UH�EH��([^_]�Z����������������SH�� H��H�I�\��H��t
H�� [�@ H�HX�S H�ك�H�� [�� ������H��X�wA���������ATUWVSH�� L�%׹ H���   H��H��H���:� 1�L�#H��f���  I�D$(H���   H�FHǃ�      ƃ�   Hǃ�      H�CH�Hǃ�      Hǃ�      Hǃ�      H�x�H�H���� H���  H���h� H���   H�VHǇ�       H���  ���   f���  ���   H�{Hǃ�      H�����  H��! H�F    H�H��(H���   �n��H���  H�� [^_]A\�H��H�� H��H��H���   �͌ H���E���L�#H��H�C    �ΐ����AUATUWVSH��(H�-u� H���   H��I��H��E���Ջ 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    �.� H��  H�H�{H��(H���   H���-o��H��H���� E��L��H��A��� W��H�H�J�H�H��t1�誥 �H��([^_]A\A]ËQ ��葥 �H��([^_]A\A]�I��H���xs��L��H�+H��H�C    H��� H��H��H���   �m�      � H���������H���א�������������AUATUWVSH��(H�-� H���   H��I��H��E���u� 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    �΢ H�o H�H�{H��(H���   H����m��H��H��袢 I�$E��H��A���U��H�H�J�H�H��t1��I� �H��([^_]A\A]ËQ ���0� �H��([^_]A\A]�I��H���r��L��H�+H��H�C    H�� H��H��H���   �� H��������H���א������������ATUWVSH�� H�-�� H���   H��H���� 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   H�C    �v� H� H�H�{H��(H���   H���ul��H��H���J� �H�� [^_]A\�H��H�$� H��H��H���   �� H������I��H����p��L��H�+H��H�C    ����������ATUWVSH�� H�BH��H�I��H�JH�P�L��H�I�PH�SH�x�I� H�H�h�H��L�H���6| H���   H��臟 H���   Hǅ�       H���   ���   f���   ���   HǇ�       ���   I�$H�{H�F    H��H�H�@�I�T$H�H�V�i��H�H�@�H���   H�� [^_]A\�I�T$H�H�R�I�L$H�H��H�C    �]����������������ATUWVSH�� H�BH��H�H��H�JH�P�H�{L��E��H�1�H�C    H�H�H�蝟 H�H��H�H�@�H�VH�       �j��H�H��H�H�H��q� E��H��H��A���oR��H�H�J�H�H��t1��� �H�� [^_]A\ËQ ���� �H�� [^_]A\�H��H����n��H��H�VH�H�R�H�NH�H��H�C    �e����ې��ATUWVSH�� H�BH��H�H��H�JH�P�H�{L��E��H�1�H�C    H�H�H�譞 H�H��H�H�@�H�VH��i��H�H��H�H�H�聞 H�U E��H��A���~Q��H�H�J�H�H��t1��(� �H�� [^_]A\ËQ ���� �H�� [^_]A\�H��H����m��H��H�VH�H�R�H�NH�H��H�C    �t����ې�UWVSH��(H�BH��H�H��H�JH�P�H�{H�1�H�C    H�H�H��ŝ H�H��H�H�@�H�VH���h��H�H��H�H�H�虝 �H��([^_]�H�VH�H�R�H�NH�H��H�C    �����H��H���1m��H���͐�����������SH�� H�� H�H��(H��H���   H�, H�AH�I�oS��H�KX�V���H�Ϡ H�KHH��H�C�>�  H��� H�C    H�H�բ H���   H��H���   辄 H��H�� [�� �SH�� H�\ H�H��(H��H���   H�� H�AH�I��R��H�KX�����H�?� H�KHH��H�C��  H�/� H�C    H�H�E� H���   H��H���   H�� [�)� ���������VSH��(H�H��H�H�@�H��H�RH�IH�T�H� H��NR��H�KX�5���H��� H�KHH��H�C��  H�FH�H�@�H�VH�H�C    H��([^Ð����������UWVSH��(H�H�p�H��H��H�H�H�X�H      ��H�H���Cx H���   H���d� H���   H���U� H���   H�MH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�W���   H�EH�UH�WH�G�Fk��H��H��([^_]Ð���������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���sw H���   H��蔙 H���   H��腙 H���   H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�W���   H�EH�UH�GH��([^_]Ð���������UWVSH��(H�iH��H��H���F� 1�H��Hǃ�       f���   H� � H�H��(H�CH�Gƃ�    Hǃ       Hǃ      H�CH�Hǃ      Hǃ      H�p�H�H��� u H���   H���q� H���   Hǆ�       H���   ���   f���   ���   Hǃ       ���   H�3 H�G    H�H��PH�CH��(H�CH��([^_]�H��H��� H��H�PH�S�� H���e��������UWVSH��(H�-�� H�qH��H��H���� 1�H�+H��f���   H�E(H��Hǃ�       ƃ�    Hǃ       Hǃ      Hǃ      Hǃ      H�CH�C    �j� H�ˬ H��H��H�CH��(H�C�L� H�= H�H��PH�CH��(H�CH��([^_]�H��H�� H��H��H�C�� H���w���H�+H��H�C    �ѐ������WVSH�� H�=�� H�qH��H��� 1�ƃ�    1�f���   H�G(H��Hǃ�       Hǃ       Hǃ      H      ǃ      Hǃ      H�;H�CH�C    �o� H�Ы 1�H��H�CH��(H�C�R� H�C H�H��PH�CH��(H�CH�� [^_�H��H�� H��H��H�C� H���~���H�;H��H�C    �ѐ�������������ATUWVSH�� H�BH��H��H�H�JH�P�M��H�I�PH�SH�x�I� H�H�h�H��L�H���6r H���   H��臕 H���   Hǅ�       H���   ���   f���   ���   HǇ�       ���   H�FI�D$    H�CH�@�H�V H�TH�H�H�@�H�V(H�H�F0H�CH�� [^_]A\Ð����WVSH�� H�BH��H�H��H�JH�P�L��H�L��H�C    H�H�H��֕ H�FH��H�CH�@�H�LH�F H�趕 H�H�H�@�H�V(H�H�F0H�CH�� [^_�H�VH�H�R�H�NH�H��H�C    ������VSH��(H�BH��H�H��H�JH�P�H�1�H�C    H�H�H��;� H�F1�H�CH�@�H�LH�F H��� H�H�H�@�H�V(H�H�F0H�CH��([^�H�VH�H�R�H�NH�H��H�C    �H�����������SH�� H�,� H�AH�Ѩ H��H�H��� H�IH�A�    H��H��| H��H�� [� �������H�� H�AH��� H��H�A�H�O� H�A�    H��H��;| �����������H�H�H�@�L�B(L�H�B0H�AH�BH�AH�@�L�B L�DH�BH�H�@�H�RH�H�A    Ð����UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���p H���   H��褒 H���   H��蕒 H���         H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�U���   H�GH�WH�EH��H��([^_]Ð������SH�� H��A��H�I�"��H��H�tHX�1�H��H�� [鰋 HX�S H�ك�H�� [陋 ���������SH�� H�H��A��H�I�h"��H��H�tHX�1�H��H�� [�]� HX�S H�ك�H�� [�F� ������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���#o H���   H���� H���   H���� H���   H�OH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�U���   H��([^_]�"��SH�� H��H�I�$��H��t
H�� [�@ H�HX�S H�ك�H�� [�V� ������H��P��,���������ATUWVSH�� L�%7� H���   H��H��H���x 1�L�#H��f���  I�D$(H���   H�Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�x�Hǃ�      H�H���l H���  H��藆 H���   H�VHǇ�       H���  ���   ���  ���   H�{Hǃ�      H�����  H� H�H��(H���   �6��H���  H�� [^_]A\�H��H�X� H��H�PH���   �Ux H�������H��L�#�֐����AUATUWVSH��(H�-�� H���   H��I��H��E���ew 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   譆 H�> H�H�{H��(H���   H���\7��H��H      ��聆 E��L��H��A���/��H�H�J�H�H��t1��)� �H��([^_]A\A]ËQ ���� �H��([^_]A\A]�H��I���;��H�+H�� H��H��H���   �w L������I����I���Ԑ�������AUATUWVSH��(H�-�� H���   H��I��H��E���%v 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   �m� H�� H�H�{H��(H���   H���6��H��H���A� I�$E��H��A������H�H�J�H�H��t1��� �H��([^_]A\A]�f.�     �Q ���ņ �H��([^_]A\A]�H��I���<:��H�+H�ғ H��H��H���   ��u L���G���I����I���Ԑ������������ATUWVSH�� H�-g� H���   H��H����t 1�H�+1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H���   �%� H��
 H�H�{H��(H���   H����4��H��H����� �H�� [^_]A\�H��H�� H��H��H���   ��t H���X���I��H���9��L��H�+��H����ATUWVSH�� H�BH�X�H�H��I��H�BL��H�H�I� H��H�h�L�H���#h H���   H���$� H���   Hǅ�       H���   ���   ���   ���   Hǃ�       ���   I�$H�^H��H�H�@�I�T$H�H�W�22��H�H�@�H���   H�� [^_]A\�I�T$H�H�R�I�L$H�H���[��������������ATUWVSH�� H�BH��H�H�H�H��H�B1�L��E��H�{H�H�      节 H�H��H�H�@�H�VH��@3��H�H��H�H�H��^� E��H��H��A�����H�H�J�H�H��t1��� �H�� [^_]A\�f.�     �Q ���� �H�� [^_]A\�H��H���^7��H��H�VH�H�R�H�NH�H���p����㐐������������ATUWVSH�� H�BH��H�H�H�H��H�B1�L��E��H�{H�H�蚁 H�H��H�H�@�H�VH��P2��H�H��H�H�H��n� H�U E��H��A�����H�H�J�H�H��t1��� �H�� [^_]A\�f�     �Q ����� �H�� [^_]A\�H��H���n6��H��H�VH�H�R�H�NH�H�������㐐������������UWVSH��(H�BH��H�H�H�H��H�BH�{1�H�H�貀 H�H��H�H�@�H�VH��h1��H�H��H�H�H�膀 �H��([^_]�H�VH�H�R�H�NH�H�������H��H���5��H���ՐSH�� H�� H�H��(H��H���   H�� H�AH�I�/��H�KP�v���H�ߌ H�K@H��H�C�^�  H�ϝ H�H�� H���   H��H���   ��p H��H�� [��� ���������SH�� H�L H�H��(H��H���   H�< H�AH�I���H�KP����H�O� H�K@H��H�C�ε  H�?� H�H�]� H���   H��H���   H�� [�Qp �VSH��(H�H��H�H�@�H��H�RH�IH�T�H�� H����H�KP�e���H�΋ H�K@H��H�C�M�  H�FH�H�@�H�VH�H��([^Ð��UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���d H���   H���      T} H���   H���E} H���   H�MH���   H���   ���   H���   ���   ���   ���   ���   ���   ���   H�W���   �4��H��H��([^_]Ð�����������SH�� H��A��H�I�+:��H��H�tHX�1�H��H�� [�Ј HX�S H�ك�H�� [鹈 ���������SH�� H�H��A��H�I��9��H��H�tHX�1�H��H�� [�}� HX�S H�ك�H�� [�f� ������UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���#c H���   H���D� H���   H���5� H���   H�OH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�U���   H��([^_]��9����������������SH�� H��H�I�<��H��t
H�� [�@ H�HX�S H�ك�H�� [�f� ������H��P�� ���������ATUWVSH�� L�%w� H���   H��H��H���l 1�L�#H��f���  I�D$(H���   H�Hǃ�      ƃ�   Hǃ�      Hǃ�      H�x�Hǃ�      Hǃ�      H�H���` H���  H���Ѓ H���   H�VHǇ�       H���  ���   f���  ���   H�{Hǃ�      H�����  H�W H�H��(H���   ��M��H���  H�� [^_]A\�H��H�P� H��H�PH���   �=l H��赼��H��L�#�֐������������AUATUWVSH��(H�-%� H���   H��I��H��E���Ek 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�            Hǃ�      H�+H���   覃 H�g H�H�{H��(H���   H���N��H��H���z� E��L��H��A���x6��H�H�J�H�H��t1��"� �H��([^_]A\A]�@ �Q ���� �H��([^_]A\A]�H��I����R��H�+H�� H��H��H���   ��j L���g���I����I���Ԑ������������AUATUWVSH��(H�-՗ H���   H��I��H��E����i 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   �V� H�  H�H�{H��(H���   H���UM��H��H���*� I�$E��H��A���'5��H�H�J�H�H��t1��у �H��([^_]A\A]� �Q ��赃 �H��([^_]A\A]�H��I���Q��H�+H��� H��H��H���   �i L������I����I���Ԑ������������ATUWVSH�� H�-�� H���   H��H���h 1�ƃ�   1�f���  H�E(H��Hǃ�      Hǃ�      Hǃ�      Hǃ�      Hǃ�      H�+H���   �� H��� H�H�{H��(H���   H���L��H��H���� �H�� [^_]A\�H��H��� H��H��H���   �h H���!���I��H���vP��L��H�+��H�������������ATUWVSH�� H�BH�X�H�H��I��H�BL��H�H�I� H��H�h�L�H����[ H���   H���4 H���   Hǅ�       H���   ���   f���   ���   Hǃ�       ���   I�$H�^H��H�H�@�I�T$H�H�W�aI��H�H�@�H���   H�� [^_]A\      �I�T$H�H�R�I�L$H�H����������������ATUWVSH�� H�BH��H�H�H�H��H�B1�L��E��H�{H�H��j H�H��H�H�@�H�VH��pJ��H�H��H�H�H��> E��H��H��A���<2��H�H�J�H�H��t1��� �H�� [^_]A\�f.�     �Q ���ŀ �H�� [^_]A\�H��H���N��H��H�VH�H�R�H�NH�H���0����㐐������������ATUWVSH�� H�BH��H�H�H�H��H�B1�L��E��H�{H�H��z~ H�H��H�H�@�H�VH��I��H�H��H�H�H��N~ H�U E��H��A���K1��H�H�J�H�H��t1��� �H�� [^_]A\�f�     �Q ���� �H�� [^_]A\�H��H���M��H��H�VH�H�R�H�NH�H���@����㐐������������UWVSH��(H�BH��H�H�H�H��H�BH�{1�H�H��} H�H��H�H�@�H�VH��H��H�H��H�H�H��f} �H��([^_]�H�VH�H�R�H�NH�H��豵��H��H���M��H���ՐSH�� H��� H�H��(H��H���   H�� H�AH�I�O3��H�KP�6���H��� H�K@H��H�C��  H�ߑ H�H��� H���   H��H���   �d H��H�� [�� ���������SH�� H�\� H�H��(H��H���   H�|� H�AH�I�2��H�KP観��H�� H�K@H��H�C莩  H�O� H�H�-� H���   H��H���   H�� [�d �VSH��(H�H��H�H�@�H��H�RH�IH�T�H��� H��>2��H�KP�%���H�� H�K@H��H�C�	      �  H�FH�H�@�H�VH�H��([^Ð��UWVSH��(H�H�p�H��H��H�H�H�X�H��H�H���CX H���   H���dz H���   H���Uz H���   H�MH���   H���   ���   H���   ���   f���   ���   f���   ���   ���   H�W���   �VK��H��H��([^_]Ð���������UWVSH��(H�=�: H��L��H���@ H��� �   H��H���� ��tH�=�: �   H����� ��uH��([^_]� H�sH���d�  E1�H��H�����  �H��([^_]�H��H���@ H���ɲ�����������UWVSH��(H�=�3 H�*L��H��H����? H��} �   H��H���� ��tH�=�3 �   H����� ��u	H��([^_]�H�sH���ä  E1�H��H���U�  �H��([^_]�H��H��� @ H���(�����������UWVSH��(H�=q9 H�*L��H��H���P? H��� �   H���� ��tH�=A9 �   H����� ��uH��([^_]� H�sH���$�  E1�H��H��趣  �H��([^_]�H��H���a? H��艱�����������UWVSH��(H�=�8 H��L��H���> H��� �   H��H���� ��tH�=�8 �   H����� ��uH��([^_]� H�sH��脣  E1�H��H����  �H��([^_]�H��H����> H���������������UWVSH��(H�=�1 H�*L��H��H���> H��{ �   H��H���� ��tH�=�1 �   H����� ��u	H��([^_]�H�sH����  E1�H��H���u�  �H��([^_]�H��H��� > H���H���
      ��������UWVSH��(H�=�7 H�*L��H��H���p= H��� �   H���� ��tH�=a7 �   H����� ��uH��([^_]� H�sH���D�  E1�H��H���֡  �H��([^_]�H��H���= H��詯�����������SH�� H�4� H��H��Y= H��H�� [�� ������������H�	� H��1= �H��� H��!= �UWVSH��(H�=1: H��L��H���= H�,� �   H��H���� ��tH�=: �   H����� ��uH��([^_]� H�sH���T�  E1�H��H����  �H��([^_]�H��H���= H��蹮�����������UWVSH��(H�=v2 H�*L��H��H��� = H��y �   H��H���� ��tH�=B2 �   H����� ��u	H��([^_]�H�sH��賠  E1�H��H���E�  �H��([^_]�H��H���= H��������������UWVSH��(H�=�8 H�*L��H��H���`< H��� �   H���� ��tH�=�8 �   H����� ��uH��([^_]� H�sH����  E1�H��H��覟  �H��([^_]�H��H���q< H���y������������UWVSH��(H�=Q8 H��L��H����; H�L� �   H��H���� ��tH�=!8 �   H����� ��uH��([^_]� H�sH���t�  E1�H��H����  �H��([^_]�H��H����; H���٬�����������UWVSH��(H�=�0 H�*L��H��H��� ; H��w �   H��H���� ��tH�=b0 �   H����� ��u	H��([^_]�H�sH���Ӟ  E1�H��H���e�  �H��(      [^_]�H��H���0; H���8�����������UWVSH��(H�=7 H�*L��H��H���: H�	� �   H���� ��tH�=�6 �   H����� ��uH��([^_]� H�sH���4�  E1�H��H���Ɲ  �H��([^_]�H��H���: H��虫�����������SH�� H��� H��H��i: H��H�� [��� ������������H�Y� H��A: �H�I� H��1: �ATUWVSH�� L�%O 1�M��L�!H��H�����A��  H�CH�k� �   H��H�H�=Y2 ��� ��tH�=I2 �   H����� ��uH�� [^_]A\�f�     H�sH���$�  E1�H��H��趜  �H�� [^_]A\�H��L�#H�����  H���$�  H���|���H��H����  H���i������������ATUWVSH�� L�%o  1�H�*M��L�!H�����A��  H�CH��� �   H��H�H�=y1 ��� ��tH�=i1 �   H����� ��uH�� [^_]A\�f�     H�sH���D�  E1�H��H���֛  �H�� [^_]A\�H��L�#H����  H���D�  H��蜩��H��H���1�  H��艩�����������ATUWVSH�� L�%�� 1�M��L�!H��H�����A�&�  H�CH��� �   H��H�H�=�0 ��� ��tH�=�0 �   H����� ��uH�� [^_]A\�f�     H�sH���d�  E1�H��H�����  �H�� [^_]A\�H��L�#H���<�  H���d�  H��輨��H��H���Q�  H��詨�����������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A�F�  H�CH��� �   H��H�H�=�/ �      ��� ��tH�=�/ �   H����� ��uH�� [^_]A\�f�     H�sH��脚  E1�H��H����  �H�� [^_]A\�H��L�#H���\�  H��脚  H���ܧ��H��H���q�  H���ɧ�����������SH�� H��� H�H��H�I��  H���=�  H��H�� [� � SH�� H��� H�H��H�I��  H��H�� [��  ��������SH�� H�t� H�H��H�I赙  H��H�� [�ؙ  ��������ATUWVSH�� L�%� 1�M��L�!H��H�����A�֘  H�CH��� �   H��H�H�=�1 ��� ��tH�=�1 �   H����� ��uH�� [^_]A\�f�     H�sH����  E1�H��H��覘  �H�� [^_]A\�H��L�#H����  H����  H���l���H��H����  H���Y������������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A���  H�CH��� �   H��H�H�=�0 ��� ��tH�=�0 �   H����� ��uH�� [^_]A\�f�     H�sH���4�  E1�H��H���Ɨ  �H�� [^_]A\�H��L�#H����  H���4�  H��茥��H��H���!�  H���y������������ATUWVSH�� L�%�� 1�M��L�!H��H�����A��  H�CH��� �   H��H�H�=0 ��� ��tH�=	0 �   H����� ��uH�� [^_]A\�f�     H�sH���T�  E1�H��H����  �H�� [^_]A\�H��L�#H���,�  H���T�  H��謤��H��H���A�  H��虤�����������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A�6�  H�CH�      �� �   H��H�H�=9/ ��� ��tH�=)/ �   H����� ��uH�� [^_]A\�f�     H�sH���t�  E1�H��H����  �H�� [^_]A\�H��L�#H���L�  H���t�  H���̣��H��H���a�  H��蹣�����������SH�� H�� H�H��H�I��  H���-�  H��H�� [�� SH�� H��� H�H��H�I�Օ  H��H�� [���  ��������SH�� H��� H�H��H�I襕  H��H�� [�ȕ  ��������SH�� H���s���H�<n H��H�H�� [Ð��������������SH�� H��蓴��H�n H��H�H�� [Ð��������������SH�� H���Ӵ��H��� H�H�� [Ð��SH�� H�t� H��H��	���H��H�� [�� ������������H�I� H������H��8H��H�
L�Q H�  I9�uH� �����@    H��8� �L$`H�D$@�L$ H��A��H�D$@H��8Ð��H��8�AoH��H�
L�Q(H��  I9�uH� �����@    H��8�H�D$@L�D$ H��)L$ A��H�D$@H��8Ð��������������HQÐ����������HQ(Ð����������H�QL�AL�IÐ��H�Q(H�Q L�A0Ð��WVSH��0H�AL�BH�q8L�AL�BH�|$(H�BH�AH�Z8L�AL�BH�BH�AL�AL�B H�BH�A L�A L�B(H�B H�A(L�A(L�B0H�B(H�A0L�A0H��H�B0H����  H��H����  H��H���ە  H��裕  �H��0[^_Ð���������1�Ð������������Hc�HQÐ�������Ð��������������Hc�HQ(Ð�������H�AH;As� �f�H�L��        H�PH�����L9�t�H�␐���H�H�`@���������L�A(L;A0��sA�H�A(�f.�     H�L�BhH��  I9�u�������    ��I�������������H�H�``���������SH�� H�d  H�H�@HH��H9�u�����H�� [�f.�     �Ѓ��t�H�S�H��H�SH�� [Ð���SH�� H�QH;QH��s�H��H�SH�� [�H�H�����H�PPH9�uH�@HH��  H9�u������� H��H�� [H��D  H���Ѓ��t�H�S�H��Ð�����������SH�� H�AH�QH��H9�sH��H�AH9�s>� H�� [�D  H�H�����H�PPH9�u=H�@HH�R  H9�uA�����H�� [�f�H�H�6  H�@HH9�t�H��H�� [H��f�H���҃��t�H�CH�S�H���Ѓ��t�H�CH�SH��H�C�j����������������SH�� H�AH;AH��sH��H�AH�� [�H�H�F���H�PPH9�u-H�@HH��  H9�t�H���Ѓ��t�H�CH�� [��     H��H�� [H�␐���AUATUWVSH��(1�M��I��I��M��~HH�=����H�-F  fD  I�T$I�D$H)�t5L��L��H)�H9�HO�I��H��E��I\$I9�hH��H��([^_]A\A]�L��I�$H�PPH9�u<H�@HH9�t�L���Ѓ��t�I�T$�H��I�T$L�KH���I9��u���� L���҃��u��H�릐��������������AUATUWVSH��(1�M��H��H��M��~8L�%]  H�N(H�F0H)�t@L��H��H)�H9�HO�I��H��D��H~(I9�H��H��([^_]A\A]�H�f�     H�H�@hL9�t��U H���Ѓ��t�H��H�      �I9��뻐������H�����H�H�@0H9�u1��f.�     H���������������H��H������A    Ð�������������H��H������A    Ð�������������H�AH9AsH�P�H�Q�@��f�     H�H��   L�@X�����I9�tމ�I�����H�AH+AuH�L��   H�R8L9�u�f�H�␐����������������Ð���������UWVSH��(H�z8H��H��H��L���S�  H�H�����H�@H9�u H��H���5�  H��H��([^_]�f�     H��H������H��H���ۏ  H��������������Ð���������L�����H�H�@L9�uH���f�     H���������������1�Ð������������H�AH9As8P�uH�P�H�Q�@��@ H�L�����L�@X�����M9�t���I���������Ð���������H�i� H�H�BH��8H��8H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A���  ���������H�� H�H��8H�A�    H�A�    H�A�    H�A�    H�A�    H�A�    �ݍ  �������������H��� H�H�BH��8H��8H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A��y�  ���������H�y� H�H��8H�A�    H�A�    H�A�    H�A�    H�A�    H�A�    �=�  �������������SH�� H�$� H�H��H�I8�Ս  H��H�� [�� ��������H��� H�H��8魍  �������������H��� H�H��8鍍  �������������SH�� H�BH�AH�BH��H��8H�I8H�A�H�B�H�A�H�B�H�A�H�B�H�A�      H�B�H�A��k�  H��H�� [Ð�H��8H��H�
L�Q H�  I9�uH� �����@    H��8� �L$`H�D$@�L$ H��A��H�D$@H��8Ð��H��8�AoH��H�
L�Q(H��  I9�uH� �����@    H��8�H�D$@L�D$ H��)L$ A��H�D$@H��8Ð��������������H�HQÐ�������H�HQ(Ð�������H�QL�AL�IÐ��H�Q(H�Q L�A0Ð��WVSH��0H�AL�BH�q8L�AL�BH�|$(H�BH�AH�Z8L�AL�BH�BH�AL�AL�B H�BH�A L�A L�B(H�B H�A(L�A(L�B0H�B(H�A0L�A0H��H�B0H����  H��H����  H��H���ۋ  H��裋  �H��0[^_Ð���������1�Ð������������Hc�H�HQÐ����Ð��������������Hc�H�HQ(Ð����H�AH;As� �f�H�L��  H�PH�����L9�t�H�␐���H�H�`@���������H�A(H;A0sf�H��H�A(����     H�L��  L�@h�����M9�t���I����H�H�``���������SH�� H�d  H�H�@HH��H9�u�����H�� [�f.�     ��f���t�H�S�H��H�SH�� [Ð��SH�� H�QH;QH��s�H��H�SH�� [�H�H�����H�PPH9�uH�@HH��  H9�u������� H��H�� [H��D  H����f���t�H�S롐��������������H��Ð�����������SH�� H�QH;QH��s.�H��H�Sf���t@H�CH;CsC� H�� [�f.�     H�H�����H�PPH9�uQH�@HH�2  H9�u-�����H�� [�f�H�H�  H�@HH9�t�H��H�� [H��f�      H����f���t�H�S�n���H�����o�����SH�� H�AH;AH��sH��H�AH�� [�H�H�F���H�PPH9�u-H�@HH��  H9�t�H����f���t�H�CH�� [��    H��H�� [H�␐���AVAUATUWVSH�� 1�M��H��I��M��~MH�-����L�%D  @ H�GH�WH9�tCH)�L��L��H��H)�H9�HN�L�4H�M���;��LwI9�lH��H�� [^_]A\A]A^� M��H�H�PPH9�uAH�@HL9�t�H����f���t�H�W�H��H�Wf���t�M�NH��fA�I9��c���뜐H������I�말���AVAUATUWVSH�� 1�M��H��I��M��~BH�-[  H�G0H�O(H9�tCH)�L��L��H��H)�H9�HN�L�4H�M���:��Lw(I9�H��H�� [^_]A\A]A^�M�H�H�@hH9�t�A�$H����f���t�H��I��I9����H�����H�H�@0H9�u1��f.�     H���������������H��H������A    Ð�������������H��H������A    Ð�������������H�AH9AsH�P��@�H�Q�f�     H�H��   L�@X�����I9�t޺��  I��H�AH�QH9�tH)�H���H�L��   H�P81�L9�t�H�␐�������Ð���������UWVSH��(H�z8H��H��H��L���c�  H�H�����H�@H9�u H��H���E�  H��H��([^_]�f�     H��H������H��H����  H��������������Ð���������L�����H�H�@L9�uH���f�     H���������������1�Ð������������H�AH9Asf9P�uH��H�A���D  H�L�����L�@X�����M9�t�      ��I���������Ð���������H��� H�H�BH��8H��8H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A��)�  ���������H��� H�H��8H�A�    H�A�    H�A�    H�A�    H�A�    H�A�    ��  �������������H�Y� H�H�BH��8H��8H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A�鉃  ���������H�	� H�H��8H�A�    H�A�    H�A�    H�A�    H�A�    H�A�    �M�  �������������SH�� H��� H�H��H�I8��  H��H�� [�� ��������H��� H�H��8齃  �������������H�i� H�H��8靃  �������������SH�� H�BH�AH�BH��H��8H�I8H�A�H�B�H�A�H�B�H�A�H�B�H�A�H�B�H�A��{�  H��H�� [Ð�UWVSH��(H�=� H��L��H���#? H�\� �   H��H���� ��tH�=� �   H����� ��uH��([^_]� H�sH���t�  E1�H��H����  �H��([^_]�H��H��H��� H��G�  H���o�  H���Ǎ���������H��H�����������UWVSH��(H�= H��L��H���c> H��� �   H��H���� ��tH�=� �   H����� ��uH��([^_]� H�sH���  E1�H��H���F  �H��([^_]�H��H��H��� H��  H���  H�������������H�������������SH�� H��� H�H��H�I�E  H���m  H��H�� [�P� SH�� H�d� H�H��H�I�  H��H�� [�8  ��������      SH�� H�4� H�H��H�I��~  H��H�� [�  ��������UWVSH��(H�=A H��L��H����> H��� �   H��H���� ��tH�= �   H����� ��uH��([^_]� H�sH���d~  E1�H��H����}  �H��([^_]�H��H��H��� H��7~  H���_~  H��跋���������H��H�����������UWVSH��(H�=� H��L��H���#> H��� �   H��H���� ��tH�=Q �   H����� ��uH��([^_]� H�sH���}  E1�H��H���6}  �H��([^_]�H��H��H��� H��w}  H���}  H��������������H�������������SH�� H��� H�H��H�I�5}  H���]}  H��H�� [�@� SH�� H��� H�H��H�I�}  H��H�� [�(}  ��������SH�� H�d� H�H��H�I��|  H��H�� [��|  ��������UWVSH��81�M��H��H�A    H����1҉AH�V� H��= H��� �   H��H�H�=e ��� ��tH�=U �   H����� ��uH��8[^_]��    H�t$(E1�H��H����{  H�T$(H���0= H���|  �H��8[^_]�H��H���S@ H��苉��H��H��� |  H���x�����������UWVSH��81�H�*M��H�A    H����1҉AH�v� H��< H��� �   H��H�H�=� ��� ��tH�=u �   H����� ��uH��8[^_]��    H�t$(E1�H��H����z  H�T$(H���P< H���8{  �H��8[^_]�H��H���s? H��諈��H��H���@{  H��蘈��      ��������UWVSH��81�M��H��H�A    H����1҉AH��� H���; H��� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]��    H�t$(E1�H��H���z  H�T$(H���p; H���Xz  �H��8[^_]�H��H���> H���ˇ��H��H���`z  H��踇����������UWVSH��81�H�*M��H�A    H����1҉AH��� H���: H�� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]��    H�t$(E1�H��H���-y  H�T$(H���: H���xy  �H��8[^_]�H��H���= H������H��H���y  H���؆����������SH�� H�T� H��H��y= H��H�� [�<� ������������H�)� H��Q= �H�� H��A= �UWVSH��81�M��H��H�A    H����1҉AH��� H��^= H�'� �   H��H�H�=% ��� ��tH�= �   H����� ��uH��8[^_]��    H�t$(E1�H��H����w  H�T$(H����< H���Hx  �H��8[^_]�H��H����? H��軅��H��H���Px  H��訅����������UWVSH��81�H�*M��H�A    H����1҉AH��� H��~< H�G� �   H��H�H�=E ��� ��tH�=5 �   H����� ��uH��8[^_]��    H�t$(E1�H��H���w  H�T$(H���< H���hw  �H��8[^_]�H��H���? H���ۄ��H��H���pw  H���Ȅ����������UWVSH��81�M��H��H�A    H����1�      �AH�� H��; H�g� �   H��H�H�=e ��� ��tH�=U �   H����� ��uH��8[^_]��    H�t$(E1�H��H���=v  H�T$(H���0; H���v  �H��8[^_]�H��H���3> H�������H��H���v  H��������������UWVSH��81�H�*M��H�A    H����1҉AH�6� H��: H��� �   H��H�H�=� ��� ��tH�=u �   H����� ��uH��8[^_]��    H�t$(E1�H��H���]u  H�T$(H���P: H���u  �H��8[^_]�H��H���S= H������H��H���u  H��������������SH�� H��� H��H��= H��H�� [�l� ������������H��� H���< �H��� H���< �1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������1�M�����AH�n� H�Ð���������SH�� H��� H��H��t  H��H�� [霺 ������������H��� H��t  �H��� H��t  �1�M�����AH�N� H�Ð���������1�M�����AH�.� H�Ð���������1�M�����AH�� H�Ð���������1�M�����AH��� H�Ð���������SH�� H�t� H��H���s  H��H�� [�̹ ������������H�I� H���s  �H�9� H��s  �1�M�����AH��� H�Ð���������1�M�����AH�>L H��H�Ð�����1�M�����AH��� H�Ð���������1�M����      �AH�n� H�Ð���������1�M�����AH��K H��H�Ð�����1�M�����AH�.� H�Ð���������SH�� H��� H��H���r  H��H�� [鼸 ������������H��� H��r  �H�y� H��r  �1�M�����AH��� H�Ð���������1�M�����AH�>K H��H�Ð�����1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������1�M�����AH��J H��H�Ð�����1�M�����AH�N� H�Ð���������SH�� H��� H��H���q  H��H�� [鬷 ������������H��� H��q  �H��� H��q  �SH�� H���C���H�\J H��H�H�� [Ð��������������SH�� H���c���H�,J H��H�H�� [Ð��������������SH�� H��裐��H��� H�H�� [Ð��SH�� H��� H��H��ِ��H��H�� [�ܶ ������������H�i� H�鱐���AVAUATUWVSH��PH��H��H���� H�����H��H� H�@ H9��}  H�FH�l$8L�D$5H��H�P�PB��H�D$8H�H�H�K�~� L�CE1�H��H��I������1�H�{ ��  �C H�H�����H�@(H9��2  H�FH�l$@L�D$6H��H�P(��A��H�D$@H�H�H�K0�� L�C0E1�H��H��I��聾��H�H�w���H�@0H9���  H�FH�l$HL�D$7H��H�P8�A��H�D$HH�H�H�K@辵 L�C@E1�H��H��I���)���H�H�����H�@H9���  H�F�@H�CHH�H�����H�@H9��U  H�F�@I�CIH���      � L�KJH��H�o@ H��H�L�B$���H�I@ H�knH�0�G8<t����   H�H�8��H�@8H9��+  H�H�CnH�FH�EH�FH�E�Ff�EH�L$HL�c�����L�s(L�k8ƃ�   ��A�����   H�L$@�������A���~_H�L$8�������A���~.H��P[^_]A\A]A^�A�$��<}������H���s���L���H�T$7H���p,���H��P[^_]A\A]A^�H�T$7H���R,���H�T$7H���B,���k���H�l$8H��H��������H���������H�l$@H��H���������H�l$HH��H��������H�����X���f�I��H��H��L�F�������E1�E1�H�D$(H�D$8H�T$5H�H���+��H�D$(H����� M��tL���d� M��tL���W� M��tL���J� �E� �H��H�D$HH�T$7H�H��}+��H��H�D$(H�D$@H�T$6H�H��b+��H�D$(�r���H���p� H���xz��H��E1��E1�E1�E1��L���H���*� �E1���2���E1�E1�����ꐐ1�H��H�A    ��H�A    �AH�~� H�1��A  H�A(    H�A0    H�A8    H�A@    f�AHƁ�    Ð��������1�H��H�A    ��H�A    �AH�� H�1��A  H�A(    H�A0    H�A8    H�A@    f�AHƁ�    Ð��������VSH��(H���"   H��H��([^��� H��H���� H���Qy���SH�� H��� ���    H��H�t*H�IH��t觱 H�K(H��t虱 H�K8H��t英 H��H�� [�k  ��������������SH�� H�D� ���    H��H�t*H�IH��t�G� H�K(H��t�9� H      �K8H��t�+� H��H�� [�>k  ��������������AVAUATUWVSH��PH��H��H��贇 H�=���H��H� H�@ H9��j  H�FL�d$8L�D$5L��H�P�<��H�D$8H�H�H�K�ް L�CE1�H��L��H���I���1�H�{ ��  �C H�H�����H�@(H9��  H�FL�l$@L�D$6L��H�P(�h���H�D$@H�H�H��������?H9�H�K0�  H��`� L�C0E1�H��L��I��蛪��H�H�����H�@0H9���  H�FL�l$HL�D$7L��H�P8�����H�D$HH�H�H��������?H9�H�K@�y  H��� L�C@E1�H��L��I���-���H�H�����H�BH9��v  H�F�@Hf�CHH�BH�����H9��F  H�F�@Jf�CJH��袁 L�KLH��H��: H��H�H�L�B$�PXH�}: L���   H��H�H�L�B�PXH�L$HH�{�����L�c(L�s8ƃ�   ��A���~sH�L$@�������A���~PH�L$8�������A���~H��P[^_]A\A]A^����<}���/���H�T$7H����&���H��P[^_]A\A]A^�H�T$7H��迢���H�T$7H��询���z���f.�     L�d$8H��L��������L�l$@H��L���������L�l$HH��L�����P���f.�     H��������fD  H����H�����E1�E1�H�D$(H�D$8H�T$5H�H��E&��H�D$(H���8� H��tH���ۭ M��tL���έ M��tcL����� �YH�D$(H�D$HH�T$7H�H�����H�D$(H�D$(H�D$@H�T$6H�H��ʡ��H�D$(�s���E1�E1�1��f���E1��H��趯 �a� H���ɱ H����t���� E1�����-���      �(���E1�E1����� �����ܐ�������1�H��H�A    ��H�A    �AH��� H��A  H�A(    H�A0    H�A8    H�A@    �AH    Ɓ�    Ð�������1�H��H�A    ��H�A    �AH��� H��A  H�A(    H�A0    H�A8    H�A@    �AH    Ɓ�    Ð�������VSH��(H���"   H��H��([^�T� H��H���I� H���s���SH�� H�$� ���    H��H�t*H�IH��t�� H�K(H��t��� H�K8H��t�� H��H�� [��e  ��������������SH�� H�Ľ ���    H��H�t*H�IH��t觫 H�K(H��t虫 H�K8H��t苫 H��H�� [�e  ��������������SH�� H���`��H��> H��H�H�� [Ð��������������SH�� H���`��H�\> H��H�H�� [Ð��������������SH�� H����`��H�� H�H�� [Ð��SH�� H�� H��H��a��H��H�� [�ܪ ������������H�ټ H���`���1�H��H�A    ��H�A    �AH�޼ H�H�A     H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    H�A`    H�Ah    H�Ap    H�Ax    Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ       Hǁ      Hǁ      Hǁ      Hǁ             Hǁ(      Hǁ0      Hǁ8      Hǁ@      HǁH      HǁP      HǁX      Hǁ`      Hǁh      Hǁp      Hǁx      Hǁ�      Ɓ�   Ð�������1�H��H�A    ��H�A    �AH�޺ H�H�A     H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    H�A`    H�Ah    H�Ap    H�Ax    Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ       Hǁ      Hǁ      Hǁ      Hǁ       Hǁ(      Hǁ0      Hǁ8      Hǁ@      HǁH      HǁP      HǁX      Hǁ`      Hǁh      Hǁp      Hǁx      Hǁ�      Ɓ�   Ð�������SH�� H��� H��H��`  H��H�� [霦 ������������H�ɸ H��`  �H��� H��`  �1�H��H�A    ��H�A    �AH��� H�H�A     H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    H�A`    H�Ah    H�Ap    H�Ax    Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�             Hǁ�       Hǁ�       Hǁ�       Hǁ       Hǁ      Hǁ      Hǁ      Hǁ       Hǁ(      Hǁ0      Hǁ8      Hǁ@      HǁH      HǁP      HǁX      Hǁ`      Hǁh      Hǁp      Hǁx      Hǁ�      Ɓ�   Ð�������1�H��H�A    ��H�A    �AH��� H�H�A     H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    H�A`    H�Ah    H�Ap    H�Ax    Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ�       Hǁ       Hǁ      Hǁ      Hǁ      Hǁ       Hǁ(      Hǁ0      Hǁ8      Hǁ@      HǁH      HǁP      HǁX      Hǁ`      Hǁh      Hǁp      Hǁx      Hǁ�      Ɓ�   Ð�������SH�� H�Ĵ H��H��i\  H��H�� [�L� ������������H��� H��A\  �H��� H��1\  �UWVSH��81�M��H��H�A    H����E1�1҉AH�� H���6��H�d� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���[  H�T$(E1�H���6��H���U[  �H��8[^_]�H��      H����9��H����h��H��H���][  H���h�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�3� H��6��H��� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���-Z  H�T$(E1�H���5��H���uZ  �H��8[^_]�H��H��� 9��H����g��H��H���}Z  H����g�������UWVSH��81�M��H��H�A    H����E1�1҉AH�S� H��;5��H��� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���MY  H�T$(E1�H����4��H���Y  �H��8[^_]�H��H��� 8��H���g��H��H���Y  H����f�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�s� H��[4��H�ı �   H��H�H�=� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���mX  H�T$(E1�H����3��H���X  �H��8[^_]�H��H���@7��H���(f��H��H���X  H���f�������SH�� H�� H��H��	7��H��H�� [�|� ������������H�� H���6���H�ٰ H���6���UWVSH��81�M��H��H�A    H����E1�1҉AH��� H���6��H�� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���=W  H�T$(E1�H���}6��H���W  �H��8[^_]�H��H����9��H����d��H��H���W  H����d�������      UWVSH��81�H�*M��H�A    H����E1�1҉AH�ӡ H��6��H�$� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���]V  H�T$(E1�H���5��H���V  �H��8[^_]�H��H����8��H���d��H��H���V  H���d�������UWVSH��81�M��H��H�A    H����E1�1҉AH�� H��+5��H�D� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���}U  H�T$(E1�H���4��H����U  �H��8[^_]�H��H���8��H���8c��H��H����U  H���%c�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�� H��K4��H�d� �   H��H�H�=2� ��� ��tH�="� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���T  H�T$(E1�H����3��H����T  �H��8[^_]�H��H���07��H���Xb��H��H����T  H���Eb�������SH�� H��� H��H���6��H��H�� [鬚 ������������H��� H���6���H�y� H���6���UWVSH��81�M��H��H�A    H����E1�1҉AH�S� H���6��H��� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���mS  H�T$(E1�H���m6��H���S  �H��8[^_]�H��H����9��H���(a��H��H���S  H���a�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�      s� H���5��H�Ĭ �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���R  H�T$(E1�H���5��H����R  �H��8[^_]�H��H����8��H���H`��H��H����R  H���5`�������UWVSH��81�M��H��H�A    H����E1�1҉AH��� H��5��H�� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���Q  H�T$(E1�H���4��H����Q  �H��8[^_]�H��H���8��H���h_��H��H����Q  H���U_�������UWVSH��81�H�*M��H�A    H����E1�1҉AH��� H��;4��H�� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H����P  H�T$(E1�H����3��H���Q  �H��8[^_]�H��H���07��H���^��H��H���Q  H���u^�������SH�� H�T� H��H���6��H��H�� [�ܖ ������������H�)� H���6���H�� H���6���UWVSH��81�M��H��H�A    H����E1�1҉AH�� H���6��H�D� �   H��H�H�=�� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���O  H�T$(E1�H���m6��H����O  �H��8[^_]�H��H����9��H���X]��H��H����O  H���E]�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�� H���5��H�d� �   H��H�H�=�� �      �� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���N  H�T$(E1�H���5��H���O  �H��8[^_]�H��H����8��H���x\��H��H���O  H���e\�������UWVSH��81�M��H��H�A    H����E1�1҉AH�3� H��5��H��� �   H��H�H�=� ��� ��tH�=�� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H����M  H�T$(E1�H���4��H���%N  �H��8[^_]�H��H���8��H���[��H��H���-N  H���[�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�S� H��;4��H��� �   H��H�H�="� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H����L  H�T$(E1�H����3��H���EM  �H��8[^_]�H��H���07��H���Z��H��H���MM  H���Z�������SH�� H��� H��H���6��H��H�� [�� ������������H�ɦ H���6���H��� H���6���AWAVAUATUWVSH��hH��H��I���Rb H�˥��H��H� H�@H9��  H�F�@!�C!H�H����H�@H9���  H�F�@"�C"H�H�q���H�@@H9���  H�F�@X�CXH�H�����H�@ H9���  H�FH�l$@L�D$<H��H�P�	��H�D$@H�H�H�K�7� L�CE1�H��H��H��袚��1�H�{ ��  �C H�H�����H�@(H9��k  H�FH�l$HL�D$=H��H�P(���H�D$HH�H�H�K0�ϑ L�C0E1�H��H��I���:���H�H����H�@0H9�       �%  H�FH�l$PL�D$>H��H�P8�I��H�D$PH�H�H�K@�w� L�C@E1�H��H��I������H�H�X���H�@8H9���  H�FL�|$XL�D$?L��H�PH����H�D$XH�H�H�KP�� L�CPE1�H��L��H��芙��H�H�Т��H�@HH9���  H�F�@\�C\H�H�����H�@PH9��2  H�F�@`�C`L���pb H�	 L�KdH��H�L�B����H�L$XH�{�����L�k(L�c8H�kH�Co��A�����   H�L$P�������A���~hH�L$H�������A���~EH�L$@�������A���~"H��h[^_]A\A]A^A_Ð���<}������H�T$?H���"����H�T$?H������H�T$?H������H�T$?H�������b���H�l$@H��H��������H�����D����H��������fD  H���������fD  H���������fD  H�l$HH��H��������H�l$PH��H���������L�|$XH��L�����)���f.�     H�����Z���1�E1�E1�H�D$(H�D$@H�T$<H�H��F��H�D$(H���9� H��tH���܎ M��tL���ώ M��tL��� H��tH��赎 谗 1�E1�H�D$(H�D$HH�T$=H�H�����H�D$(�{����n���H���� H����U����1�E1�E1��1�E1�E1�1��K���H��衐 �1�H�D$(H�D$PH�T$>H�H����H�D$(�1�E1�������1���H��H�D$XH�T$?H�H��X��H���H��1���1���C������1�H��H�A    ��H�A    �AH�� H�1�f�A �A" H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �A!      o Ð������������1�H��H�A    ��H�A    �AH��� H�1�f�A �A" H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Ao Ð������������VSH��(H���"   H��H��([^�� H��H���ٌ H���AT���SH�� H�� �yo H��H�t8H�IH��t蚌 H�K(H��t茌 H�K8H��t�~� H�KHH��t�p� H��H�� [�F  ���SH�� H��� �yo H��H�t8H�IH��t�:� H�K(H��t�,� H�K8H��t�� H�KHH��t�� H��H�� [�#F  ���AWAVAUATUWVSH��hH��H��I����[ H�;���H��H� H�@H9��  H�F�@!�C!H�H�����H�@H9���  H�F�@"�C"H�H����H�@@H9���  H�F�@X�CXH�H����H�@ H9���  H�FH�l$@L�D$<H��H�P�9��H�D$@H�H�H�K�g� L�CE1�H��H��H���ғ��1�H�{ ��  �C H�H�(���H�@(H9��k  H�FH�l$HL�D$=H��H�P(����H�D$HH�H�H�K0��� L�C0E1�H��H��I���j���H�H�P���H�@0H9��%  H�FH�l$PL�D$>H��H�P8�y��H�D$PH�H�H�K@觊 L�C@E1�H��H��I������H�H�Ƞ��H�@8H9���  H�FL�|$XL�D$?L��H�PH�!��H�D$XH�H�H�KP�O� L�CPE1�H��L��H��躒��H�H�@���H�@HH9���  H�F�@\�C\H�H����H�@PH9��2  H�F�@`�C`L���[ H�9 L�KdH��H�L�B�F���H�L$XH�{�����L�k(L�c8H�kH�Co"      ��A�����   H�L$P�������A���~hH�L$H�������A���~EH�L$@�������A���~"H��h[^_]A\A]A^A_Ð���<}������H�T$?H���R����H�T$?H���B���H�T$?H���2���H�T$?H���"���b���H�l$@H��H��������H�����D����H��������fD  H���������fD  H���������fD  H�l$HH��H��������H�l$PH��H���������L�|$XH��L�����)���f.�     H�����Z���1�E1�E1�H�D$(H�D$@H�T$<H�H��v ��H�D$(H���i� H��tH���� M��tL����� M��tL���� H��tH���� ��� 1�E1�H�D$(H�D$HH�T$=H�H�� ��H�D$(�{����n���H���� H���$O����1�E1�E1��1�E1�E1�1��K���H���щ �1�H�D$(H�D$PH�T$>H�H�����H�D$(�1�E1�������1���H��H�D$XH�T$?H�H�����H���H��1���1���C������1�H��H�A    ��H�A    �AH�n� H�1�f�A �A" H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Ao Ð������������1�H��H�A    ��H�A    �AH�� H�1�f�A �A" H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Ao Ð������������VSH��(H���"   H��H��([^�� H��H���	� H���qM���SH�� H�T� �yo H��H�t8H�IH��t�ʅ H�K(H��t輅 H�K8H��t讅 H�KHH��t蠅 H��H�� [�?  ���#      SH�� H��� �yo H��H�t8H�IH��t�j� H�K(H��t�\� H�K8H��t�N� H�KHH��t�@� H��H�� [�S?  ���AWAVAUATUWVSH��hH��H��H���rU H�����H��H� H�@H9��8  H�F�@"f�C"H�H����H�@H9��5  H�F�@$f�C$H�H�O���H�@@H9��  H�F�@X�CXH�H�~���H�@ H9��  H�FL�d$@L�D$<L��H�P�g��H�D$@H�H�H�K蕄 L�CE1�H��L��H��� ���1�H�{ �(  �C H�H�����H�@(H9���  H�FL�l$HL�D$=L��H�P(����H�D$HH�H�H��������?H9�H�K0��  H��� L�C0E1�H��L��I���R~��H�H�����H�@0H9��O  H�FL�l$PL�D$>L��H�P8豌��H�D$PH�H�H��������?H9�H�K@�r  H�詃 L�C@E1�H��L��I����}��H�H�
���H�@8H9��  H�FL�l$XL�D$?L��H�PH�C���H�D$XH�H�H��������?H9�H�KP��  H��;� L�CPE1�H��L��I���v}��H�H�l���H�@HH9���  H�F�@\�C\H�H�;���H�@PH9��n  H�F�@`�C`H����T H�% L�KdH��L�H�L�BA�RXH�L$XH�{�����L�c(L�s8L�{H�Cz��A�����   H�L$P�������A���~gH�L$H�������A���~DH�L$@�������A���~!H��h[^_]A\A]A^A_����<}�������H�T$?H���=�����H�T$?H���v���H�T$?H���v���H�T$?H����u���c����     H���������fD  H���������fD  H�������$      ��fD  L�d$@H��L��������L�l$HH��L�����]���L�l$PH��L��������f.�     H��������fD  L�l$XH��L���������H�����L���E1�E1�E1�H�D$(H�D$@H�T$<H�H��S���H�D$(H���F� H��tH���� M��tL���܀ M��tL���π M��tL��� 轉 H�D$(H�D$XH�T$?H�H���t��H�D$(H�D$(H�D$PH�T$>H�H���t��H�D$(H�D$(H�D$HH�T$=H�H��t��H�D$(�F���H���Ʉ H����G��E1���� ��E1�E1�E1���� ���
���E1�E1�E1�1����������E1��q������ډ E1�E1��|���E1�E1��T�������H���8� �!����������������������1�H��H�A    ��H�A    �AH�>� H��A  �A"    H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Az Ð�����������1�H��H�A    ��H�A    �AH��� H��A  �A"    H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Az Ð�����������VSH��(H���"   H��H��([^��~ H��H���~ H���!F���SH�� H�$� �yz H��H�t8H�IH��t�z~ H�K(H��t�l~ H�K8H��t�^~ H�KHH��t�P~ H��H�� [�c8  ���SH�� H�Ē �yz H��H�t8H�IH��t�~ H�K(H��t�~ H�K8H��t��} H�KHH��t��} H��H�� [�8  ���AWAVAUATUWVSH��hH��H��H���N H�����H��H� H�@H9��8  H�F�@"%      f�C"H�H����H�@H9��5  H�F�@$f�C$H�H�?���H�@@H9��  H�F�@X�CXH�H�n���H�@ H9��  H�FL�d$@L�D$<L��H�P�	��H�D$@H�H�H�K�E} L�CE1�H��L��H��谅��1�H�{ �(  �C H�H�����H�@(H9���  H�FL�l$HL�D$=L��H�P(�υ��H�D$HH�H�H��������?H9�H�K0��  H���| L�C0E1�H��L��I���w��H�H�����H�@0H9��O  H�FL�l$PL�D$>L��H�P8�a���H�D$PH�H�H��������?H9�H�K@�r  H��Y| L�C@E1�H��L��I���v��H�H�����H�@8H9��  H�FL�l$XL�D$?L��H�PH����H�D$XH�H�H��������?H9�H�KP��  H���{ L�CPE1�H��L��I���&v��H�H�\���H�@HH9���  H�F�@\�C\H�H�+���H�@PH9��n  H�F�@`�C`H���M H�� L�KdH��L�H�L�BA�RXH�L$XH�{�����L�c(L�s8L�{H�Cz��A�����   H�L$P�������A���~gH�L$H�������A���~DH�L$@�������A���~!H��h[^_]A\A]A^A_����<}�������H�T$?H���������H�T$?H����n���H�T$?H���n���H�T$?H���n���c����     H���������fD  H���������fD  H���������fD  L�d$@H��L��������L�l$HH��L�����]���L�l$PH��L��������f.�     H��������fD  L�l$XH��L���������H�����L���E1�E1�E1�H�D$(H�D$@H�T$<H�H�����H�D$(H����{&       H��tH���y M��tL���y M��tL���y M��tL���ry �m� H�D$(H�D$XH�T$?H�H��m��H�D$(H�D$(H�D$PH�T$>H�H��xm��H�D$(H�D$(H�D$HH�T$=H�H��[m��H�D$(�F���H���y} H���@��E1���ǂ ��E1�E1�E1��赂 ���
���E1�E1�E1�1����������E1��q�����节 E1�E1��|���E1�E1��T�������H����z �!����������������������1�H��H�A    ��H�A    �AH�� H��A  �A"    H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Az Ð�����������1�H��H�A    ��H�A    �AH��� H��A  �A"    H�A(    H�A0    H�A8    H�A@    H�AH    H�AP    H�AX    �A`    �Az Ð�����������VSH��(H���"   H��H��([^�tw H��H���iw H����>���SH�� H�� �yz H��H�t8H�IH��t�*w H�K(H��t�w H�K8H��t�w H�KHH��t� w H��H�� [�1  ���SH�� H��� �yz H��H�t8H�IH��t��v H�K(H��t�v H�K8H��t�v H�KHH��t�v H��H�� [�0  ���SH�� H�$� H��H��0  H��H�� [�|v ������������H��� H��q0  �SH�� H�D� H��H��Y0  H��H�� [�<v ������������H�� H��10  �SH�� H��� H��H��i�  H��H�� [��u ������������H�i� H��A�  �SH�� H��� H��H��8��H��H�� [�'      �u ������������H��� H��8���SH�� H�$� H��H��/  H��H�� [�|u ������������H��� H��q/  �SH�� H�D� H��H��Y/  H��H�� [�<u ������������H�� H��1/  �SH�� H�� H��H��i�  H��H�� [��t ������������H�� H��A�  �SH�� H�4� H��H��)�  �   H��H�� [��t �������H�	� H���  �SH�� H�$� H��H��.  H��H�� [�|t ������������H��� H��q.  �SH�� H�D� H��H��Y.  H��H�� [�<t ������������H�� H��1.  �SH�� H�� H��H��i�  H��H�� [��s ������������H��� H��A�  ���s �����������Ð��������������H�ɜ Ð�������H�ɜ Ð�������AWAVAUATUWVSH��(�AH��$�   H��$�   %�   L��M��I����H)�� ��   ����   H�t H��u]M��ujH��([^_]A\A]A^A_É�D  A8Fiu�H��~�A�UA:��   ��  A���   8���  H�t H��t�     I�؉�H���C���M��t�M��L��H��H��([^_]A\A]A^A_�0���H��u+H���j���H�L5 I�؉�H��([^_]A\A]A^A_����� I��L��H�������H���1������    H���   �4D �x8 I��t+A�E A8Fft
A8Fd�����E L�f�H��I�������f�L�=����H���A���I�L�@0�-   M9���   A�U 8�t�A�~8 ��   L������I�L�@0�+   M9���   A�U 8�t�A�~8 ����(      �L�������I�L�@0�0   M9���   A8E �I���H���?���A�~8 �g����x   L���~���A�U8�tEA�~8 �X����X   L���]���A�U�I��� �+   L��A���e����-   L��A���$���A�E L�f�H��I���E�A�E��E������0   L��A���U�����������������AVAUATUWVSH��0�AH��$�   H��$�   %�   L�ǉ�I��H)�� �&  L�$��t2J�'H��t1�f�f�4GH��H9�u�M����   H��0[^_]A\A]A^�H���   L�L$(�B �-   I��H� L���PPL�L$(fA9�  I��+   L���PPL�L$(fA9��   I�L�L$(�0   L���PPL�L$(fA9�^���H���T���I��x   L���PPL�L$(fA9A��   I�L�L$(�X   L���PPL�L$(fA9A��   J�'H������O�D- L��H��0[^_]A\A]A^�����     L�d- H��u9L�1�H��������     f�4GH��H9������f�4GH��H9�u������H��M��L������L�1�H��u�����f�L�m�H��I���o���A�L�m�H��I��f�G�A�A�f�G��M�������������H�ɒ Ð�������W1�M��I��H�A     ��H�A(    �AH�� H��H��H���A!�H��H��� D�AHD�1�H�Q0H�Q9�    H���H�I��9  �    A�B8 H���H�AƂ9   _Ð�W1�H�|$0 ��H��H�A     �AH� H�A(    H��M��H���A!�M��H��� D�ILD�1�L�A0L�A9�    L���H�L��9  �    �B8 L���H�Ƃ9   _ÐSH�� H���   H��)      H�� [��m ������SH�� H�� H��H�H�I�'  �{ tH�K0H��t�m H��H�� [�'  ����WVSH�� 1�H���f��DH��H���   to���HJ�����u��F 1ۉ��V;��f��^�   H��H��   u�1ۿ   f.�     �ى���H��f��^�  �
���f��^�  H��H��u�H�� [^_��F뛐���������SH�� 1�M��H��H�T$8���AH�Q� H�H�L$8�$&  �C H��H�C�$����H�� [Ð������������VSH��(1�H��H�����AH�� H��%  H��H�C�C H��([^�����H��H��� H��H�PH��N&  H���3��������SH�� H��� H��H�H�I��%  H��� H��H��H��&  H��H�� [��k ��SH�� H�t� H��H�H�I�%  H�n� H��H��H�H�� [��%  ����������SH�� H��� H�M   �X��H�a� H�; tH�� [�D  H�Y� �   ��  H�x� H�A� H�H�H�� [Ð����H��(H�%� �   �  H�� H�� H�H�3� H�H��(Ð����������H��(��t��?u��w"H� �ɋ���H��(�������u���H��(�H��� �@ ����������������AWAVAUATUWVSH��(H�� L�2L�j���    L�bH��H��� H��H��1�L�5�� H��� �^�  ���� H�o� H�{�����H�o� H��H�D� ���    H��H�o� �j#  H�s� ��c� H�t� H�{����H�D� E1�H��H��� H��� 1����    L�-�� H��*      H��� ��������� H�=� H�{�T���H�m� E1�H��H�?� H�x� 1��t�    L�%u� H��H�Z� �E����U� H��� H�{�����H�6� H��H�K� �ɚ    H��H��� ���� H��� H�{����H��� H��H�,� ���    H��H��� ���� H��� H�{����H�x� H��H�]� �+�    H��H�� ��� H��� H�{�@���H��� H��H�n� �   �$�  ��d� H�e� H�{����H�E� H��H��� H��� 1����    H�nH�~ H�v(H��H�p� H�-y� ��  ��d� H�5� L�{����H�E� I��H�
� �X�    H��H�E� � !  H�I� ��9� H�:� L�{�a���H�� E1�I��H�\� H��� 1����    H�=�� H��H��� ������� H�� L�{�
���H�c� E1�I��H�� H�n� 1��j�    H�5k� H��H�P� �����K� H��� L�{����H�,� I��H�� ���    H��H�|� ��|� H�m� L�{�t���H�]� I��H��� �p�    H��H�]� ��]� H�N� L�{�5���H�>� I��H�#� ��    H��H�ޗ ��ޗ H��� L�{�����H��� �   I��H�?� ��  ��:� H�+� L�{�����H�+� H�� I��L�{����H��� M�4�L�s����H�|� M�,�L�k���+      �H��� M�d� L�c�j���H�c� I�,�H�k�V���H�_� H�[H�|� �A���H�4�H��([^_]A\A]A^A_�H��� H���  H����,��H��� H���v  H����,��H�W� H���_  H���,��H��� H���H  H���,��H�i� H���1  H���,��H�� H���  H���r,��H��� H���  H���[,��H�$� H����  H���D,������AWAVAUATUWVSH��8L��$�   H�˹   H��M��L����d H�H���@    H��� H�G    H��H��H��g�  ��GH�{� L�s�����   I�<�L�t$(�d L��H��H��G    H�D$(H�3� H��H��  H�G��GH�w� L�{�����   I�<��@d H�E1�H���@    H�y� H�G    H��H��H��������GH�F� L�{�]����   I�<���c H�E1�H���@    H�8� H�G    H��H��H��Q�����GH�� L�{�����   I�<��c H���@    H�M� H��H���GH��� L�{������   I�<��cc H���@    H�2� H��H���GH��� L�{�����   I�<��(c H���@    H�g� H��H���GH��� L�{�[����    I�<���b H�E1�I��H��H�����  ��GH�}� L�{�$����   I�<��b H�H���@    H��� H�G    H��H��H����  ��GH�_� L�{������   I�<��hb L��H��H��G    H�D$(H�� H��H��p  H�G��GH�`� L�s���,      ��   I�<��b I�U M��H���@    H�q� H�G    H��H��H��:�����GH�>� L�s�5����   I�<���a I�U M��H���@    H�/� H�G    H��H��H������GH��� L�c������   I�<��ua H���@    H�4� H��H���GH��� L�c�����   I�<��:a H���@    H�� H��H���GH��� L�c�m����   I�<���` H���@    H�N� H��H���GH��� L�c�2����    I�<���` H�E1�I��H��H����  ��GH�d� H�[�����H�<�H��8[^_]A\A]A^A_�H��H���K  H���3` H���'��H��H��� ` H���'�������������Ɛ�����������WVSH��0��u ��H��H��L����   H��� H�L$(�0������Z  H��� H�
H��u#�w�    �K���H9���   H��H�
H��tV�1���H9�H�Ju��#���H�WH��H�<� ��   H��t	H�H���PH�L$(�Y�������   H��0[^_�f�     H�GH�<� u���FH�GH�4���fD  H��t �Te ���+���H�Ş 1��N���H��t �f H�j �Vu��� ����H�
�x���H�WH��H��H�<� �R���H�F�� H�WH���H�4��F����� H�GH�4��5���H�=�M �   ��_ L�PB��H�8H�V H���g H�=M �   �_ L��A��H�8H�� H���g H��H��u,�6a H��s H���c H���%��H�L$(H���b,��H���z%������������AWAVAUATUWVSH��(-      M��H��L���  H���y���H��H�FH��H9���   L�cL�nH��������N�<�    I9�H������LG�L���] H�NH��H��tL�F1� I��H��H��H9�u�I9�vH��H�T� �H�     H��H9�u�L��L�v�d] L�FM��tL�N1�D  I��H��H��L9�u�M9�vJ��H�L� �H�    H��H9�u�M��L�fH�~H�FtL����\ M��tL����\ ��EH�FH�<�H�H����   H��� H�
H��u$�oH�J�G���H9���   H��H�
H����   �)���H9�u�H�JL�F����I��H�; ��   H�RH������I����@H���i��   L�#H���htzH�~ H�/tP1�H�F��     H�FH�8    H��H9^v*H��H�<�    H��t���iu�H��P��f.�     H��([^_]A\A]A^A_�H��f.�     H�H���RH�~ H�/�y������    H�
L�F�4���I��H�; t�H�H�������I����@H���i�"���H��P����H��P����H���] �_ ����H���y] H���![ �d H���d] �_ �����H���R] �m_ �����H���@] �[_ ����H��H��u��] H���@_ H���H"�������ܐ�H��(I��L��M���^���H�JH��H9�rH�RL��M��tL��L��H��(����H��� �� ���������WVSH�� L��M� H��H��M��t�     H��H��H������L�M��u�H�� [^_ÐATUWVSH�� H�BH��H�AH��������H��H9�D�H�A    H�A    H�A     H��    .      H������HG��Z L�CH�CM��L��tO1��@ H�CH�OH��H��H��t	��AL�CH��I9�w�H��������J��    I9�H������HG��Y H�{ H�Ct-1��	D  H�CH�OH��H��H��t��AH��H9Swܹ0   �bY H�C H�P0f.�     H�     H��H9�u�1�H�G H�0H��t>����L�c H�hH��I��Y I�$H�C I��H�0H�G H�0H���I���H��0u�H�� [^_]A\�H��� [ H���  �a H���] H��� �����AWAVAUATUWVSH��X�H��H�A.   H�� H��p  H��f�H�     H��H9�u�H�KH�u} H��p  H��H�     H��H9�u�H�KH�} H�Q0H��f�     H�     H��H9�u�H�K H��w H��| �)  A�   E1�1�� H��w f�]w �����H��� L�jw H�������H�[~ �   �q�  H��� L�C~ H������H��� 1�1��ip  L�5Bp f��p H��m �2p    H�/p     H��H�(p     H�	p H�"� H�p     H�p     H�p     H��H�p     �Sp  �im    H�Zm L�5cm 莠  H��� L�@m H�������H��� L�z H���u    H�6� H��H�[ ����H��� L�h H���c    H�$� H��H�I �t���H�-� �K}    H��H�8} �  H��� L�%} H��H�+} �6���H�� 1�E1���s  L�-�s f��s 1�H�,n ��s    H�/      �s     H��H��s     H�as H�Z� H�ws     H�ts     H�qs     H��H�js     H�gs     H�ds     H�as     �_s     �gs  ��m    H��m L�-�m �+  H�t� L�mm H���E���H��� L�%7s E1�1�H�km �)s    H�&s     H�#s     H���"s  H��r 1�f�s H�y� H�s     H�s     H� s     H��H��r     H��r     H��r     H��r     ��r     ��r  ��l    H��l L�%�l ��  H��� L��l H���T���H�m� L�Fk H���Ak    H�� H��H�'k �"���H�[� L�4k H���/k    H� � H��H�k �����H�� A�   �!n    H�n H�n     H� k H�n     H�
n     H�n     H��H��m H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     H��m     0      H��m     H��m     H��m     H��m     H��m     H�~m     H�{m     �|m  �O���H�h� L��h H������H��� L�+h H���&h    H�7� H��H�h �g���H�� L�h H���h    H��� H��H��g �5���H�Ng �   �t�  H��� L�6g H������H��r �   �m���H��� L��r H�������H��w �   趦  H�� L��w H�������H��� H�-j 1��j    H�g �j  H��i     H��i     H��H��i     H��i H�U� H��i     H��i     H��i     H����i     �Wj  ��f    H��f H�-�f �B�  H��� L��f H�������H�%� L��x H����x    H�j� H��H��x �����H�� L��x H����x    H�X� H��H�}x ����H�a� ��v    H��H�|v �  H��� L�iv H��H�ov �Z���H��� H�=�m E1�1�H��g ��m    H��m     H��m     H����m  H��m H��� ��m     H��m     H��m     H��H��m     H��m     H��m     H��m     H��m     ��m     ��m  ��f    H��f H�=�f ��  H��� L��f H���h���H��� H�5Zm E1�1�H��f �Lm    H�Im     H�Fm     H���Cm  H�m H��� �-m1           H�(m     H�%m     H��H�m     H�m     H�m     H�m     H�m     �m     �#m  �'f    H�f H�5!f �  H��� L��e H���v���H��� L�xd H���sd    H�D� H��H�Yd �D���H��� L�fd H���ad    H�2� H��H�Gd ����H�K� A�   ��h    H��h H��h     H�bd H��h     H��h     H��h     H��H��h H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H��h     H�h     H�|h     H�yh     H�vh     H�sh     H�ph     H�mh     H�jh     H�gh     H�dh     H�ah     H�^h     H�[h     H�Xh     H�Uh     H�Rh     H�Oh     H�Lh     H�Ih     H�Fh     H�Ch     H�@h     H�=h     �>h  �����H��� L�Cb H������H��� L�]a H���Xa    H�i� H��H�>a ����H�B� L�Ka H���Fa    H��� H��H�,a �W���H��` �   �f�  H��� L�x` H���0���H�� L�a H����` 2         H�>� H��H��` �����H��� L��` H����`    H��� H��H��` �����H�T$ H��L�t$ L�l$(L�d$0H�l$8H�|$@H�t$H�����H�:� L�{�1���H��� M�4�L�s����H��� M�,�L�k�	���H�"� M�d� L�c�����H��c I��H��� L�c�ٴ��H�r� I�,�H�k�Ŵ��H�n� H�|� H�{谴��H��� H�[H�4�H�5�d 蕴��H�4�H��X[^_]A\A]A^A_�H��H���H�Qa H��H����  H��H����   �K H��` H��H���  ��H��` H��H���  ��H��o H��H���  �H��` H��H���v  �H��^ H��H���b  �H�)o H��H���N  �s���H��^ H��H���7  �\�������������������VSH��(H�AH��H��tKH�y t<1�� H�CH��H9sv"H��H��t���iu�H��P��f.�     H��tH���G H�CH��tGH�{ t81��H�CH��H9sv!H��H��t���iu�H��P��f�     H��tH���SG H�C 1�H��t8�     H�0H��t	�2G H�C H��H��0u�H��tH��H��([^�G �H��([^�H���QI �lK �h���H���?I �ZK ����H��H��u��I ���P������������������H�Y� Ð�������H��(H�u   H�~z �i���H�bz H��(Ð������������1�Ð������������WVH��(H�=� H�    H�ֹ   ��� ��uH��(^_�H�ӟ ��  ������H��� E1�H��y ��������������3      H�    Ð�������1�Ð��������������E �����������Ð��������������UWVSH��XH��H���������H��H�D$(��������   H��� H�H�(��H�H�\$0H�H��H���\���H�� H���=�����u9H�L$0H��H9�t�fE H�L$(�\�����u+H��H���   H��H��X[^_]ÐH�T$01��t�����},��H�=&4 �   �|F L��(��H�8H��� H���CN H�L$(H���F��H���^��H��H��u���G ����������������H��(����H��� H�yi H��   H�ji H��(Ð����H�Ð�����������H�H��� Ð����WVSH�� H�    H������H�5s� H�,� H�H�H;t5�<��H��H��������uWH��� H�H��H��(�����uH�� [^_��� H�� [^_ù   �fE H��2 H�L��'��H��H��� �&M �1+��H��H��u��F ���<��������������SH�� H���+tH�� [�H������H��H�� [�C �������SH�� H��H�
��H���+tH�H�H�� [�H��H�T$8H�D$0�J���H���RC H�T$8H�D$0H�H�H�� [Ð�����������SH�� H�AH��H����   �@!.H�C�@",H�SH��� H�BH�SH�B    H�SH�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�� H�S� �B\H�S�B`H��� L� 1�f.�     A� H�S�LdH��H��u�H�� [� �p   �B H��� �@    H�@    H�@    H�Q�@" H�1�f�P4       H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@o H�C����������������VSH��(1�M��H�QH����E1�1҉AH�; H��t����H��([^�H��H������H���������������VSH��(1�M��H�A    H�����AH��: H��%����H��([^�H��H���R���H���������������VSH��(1�H��H�A    H����E1�1҉AH�x: H�������H��([^�H��H�������H���U�������VSH��(1�M��H�QH����E1�1҉AH�,: H������H��([^�H��H������H���	�����������VSH��(1�M��H�A    H�����AH��9 H��5����H��([^�H��H���b���H���������������VSH��(1�H��H�A    H����E1�1҉AH��9 H�������H��([^�H��H������H���e�������VSH��(H���"   H��H��([^��? H��H����? H���1���VSH��(H�3� H��H��H�H�IH��tH��PH��H��([^����H��H������H���������������SH�� H�AH��H����   �@!.H�C�@",H�SH�ԁ H�BH�SH�B    H�SH�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�F� H�S� �B\H�S�B`H�?� L� 1�f.�     A� H�S�LdH��H��u�H�� [� �p   ��> H��� �@    H�@    H�@    H�Q�@" H�1�f�P H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X   5       �@`    �@o H�C����������������VSH��(1�M��H�QH����E1�1҉AH��7 H��t����H��([^�H��H�������H���9�����������VSH��(1�M��H�A    H�����AH�}7 H��%����H��([^�H��H������H����������������VSH��(1�H��H�A    H����E1�1҉AH�(7 H�������H��([^�H��H���=���H����������VSH��(1�M��H�QH����E1�1҉AH��6 H������H��([^�H��H�������H���I�����������VSH��(1�M��H�A    H�����AH��6 H��5����H��([^�H��H������H����������������VSH��(1�H��H�A    H����E1�1҉AH�86 H�������H��([^�H��H���M���H����������VSH��(H���"   H��H��([^�< H��H���	< H���q���VSH��(H��� H��H��H�H�IH��tH��PH��H��([^�����H��H�������H���)�����������SH�� H�AH��H����   �.   �,   f�P"H�Cf�H$H�CH�
~ H�HH�CH�@    H�SH��} H�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H�u� H�S� �B\H�S�B`H�n� L� 1�f�     fA� H�Sf�LBdH��H��u�H�� [Ð��   �; H�/� �@    H�@    H�@    H�Q�@  H��@"    H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@z H�C��������������VSH��(1�6      M��H�QH����E1�1҉AH�l4 H��d����H��([^�H��H������H���i�����������VSH��(1�M��H�A    H�����AH�4 H������H��([^�H��H�������H���������������VSH��(1�H��H�A    H����E1�1҉AH��3 H�������H��([^�H��H���m���H���� �������VSH��(1�M��H�QH����E1�1҉AH�|3 H��t����H��([^�H��H���!���H���y �����������VSH��(1�M��H�A    H�����AH�-3 H��%����H��([^�H��H�������H���* ������������VSH��(1�H��H�A    H����E1�1҉AH��2 H�������H��([^�H��H���}���H������������VSH��(H���"   H��H��([^�D8 H��H���98 H�������VSH��(H��� H��H��H�H�IH��tH��PH��H��([^����H��H������H���Y������������SH�� H�AH��H����   �.   �,   f�P"H�Cf�H$H�CH�:z H�HH�CH�@    H�SH�!z H�B(H�SH�B0    H�SH�B8H�SH�B@    H�SH�BHH�CH�@P    H�C�@X    H��� H�S� �B\H�S�B`H��� L� 1�f�     fA� H�Sf�LBdH��H��u�H�� [Ð��   �67 H�o� �@    H�@    H�@    H�Q�@  H��@"    H�@(    H�@0    H�@8    H�@@    H�@H    H�@P    H�@X    �@`    �@z H�C��������������VSH��(1�M��H�QH����E1�1҉AH�1 H��d����H��7      ([^�H��H���A���H���������������VSH��(1�M��H�A    H�����AH��0 H������H��([^�H��H�������H���J�������������VSH��(1�H��H�A    H����E1�1҉AH�h0 H�������H��([^�H��H������H������������VSH��(1�M��H�QH����E1�1҉AH�0 H��t����H��([^�H��H���Q���H���������������VSH��(1�M��H�A    H�����AH��/ H��%����H��([^�H��H������H���Z�������������VSH��(1�H��H�A    H����E1�1҉AH�x/ H�������H��([^�H��H������H�����������VSH��(H���"   H��H��([^�t4 H��H���i4 H��������VSH��(H�� H��H��H�H�IH��tH��PH��H��([^�<���H��H���1���H���������������H�	�4 ��������H�H�AH9�tH����3 Ð����������AWAVAUATUWVSH��8H��������H��$�   H��H�IL�L��H)�H9��V  H�I��M)�L�CJ�,)L9���  L�CI9��N  L�4I��H�I)�A��H9���A!�L9�voE��t*I�6I��I�>�9  M��L��$�   蠢��L��$�   H��tH���  I��L��L��胢��H�H�k�( H��H��8[^_]A\A]A^A_�@ H�I9�w�H����   H9���   H����   L��I��L��L��$�   ����E��L��$�   t�f�     I�6I��I�>��   M��L��$�   ����L��$�   H9��Z���I�9L�H9���   L9���   K�)H���� 8        I��L��諡���#���fD  H�|$ I��H����  ����A�A�������������D  A�   �n���D  A�A�E���j����;���H��t�I��L��L���/�������f����@���fD  L)�H��t:H��tI��L��L�������I�>I��I�6I)�I��tM���d��������Z���A�A������G����A��<���H�Ȃ ���  �������H)�H������@H��   �M�ÐH�QÐ����������H�Ð�����������H�Ð�����������H�Ð�����������H�Ð�����������VSH��(H��D��H��H�T$HI��w6H�M��tI��tH@��H�������L�D$HH�L�CB�  H��([^�@ H�T$HE1���  L�D$HH�L�C�D  @�0L�D$HH�L�CB�  H��([^Ð����WVSH��0L��H��H��H)�H��H�\$(wBH��H�u��H�\$(H�H�^� H��0[^_�H��u0H�^� H��0[^_��    H�T$(E1��#  H�T$(H�H�VI��H��H���)���H�\$(H�H�^� H��0[^_ÐWVSH��0L��H��H��H)�H��H�\$(wBH��H�u��H�\$(H�H�^� H��0[^_�H��u0H�^� H��0[^_��    H�T$(E1��  H�T$(H�H�VI��H��H��艞��H�\$(H�H�^� H��0[^_ÐWVSH��0H��H��H��u	M����   L��H)�H��H�\$(wDH��H�u��H�\$(H�H�^� H��0[^_�H��u5H�^� H��0[^_�f�     H�T$(E1�H����  H�T$(H�H�VI��H��H���֝��H�\$(H�H�^� H��0[^9      _�H�7� ���  ��WVSH��0H��H��H��u	M����   L��H)�H��H�\$(wDH��H�u��H�\$(H�H�^� H��0[^_�H��u5H�^� H��0[^_�f�     H�T$(E1�H���  H�T$(H�H�VI��H��H������H�\$(H�H�^� H��0[^_�H�w ��  ��H�AÐ����������H�H�Q� Ð���I)�I��tM��uÐ黜����Ð����I)�I��tM��uÐ雜����Ð����I)�I��tM��uÐ�{�����Ð����I)�I��tM��uÐ�[�����Ð����H��(H�AH9t#H�AH9Ar	H��(�@ 1��9  �H��(� �   ��H����. �H��(��0 �������ATUWVSH��0H����������$�   L��L�IL�H��H��L)�H9���   H�	H�CI��M)�M�H9���   H�CL9�rgI�(I)�t$I9�tH�J�H�I����   M���u���H�H��tH�H��t\@��I���P���H�H��L�cB�! H��0[^_]A\�fD  E1�H��H�t$ H���  H��H�t�� �   �j���fD  @�9H���     �H���H�t��y���H��| ��  ��H��Ð�����������E�������������H��(L�AL9�sH�H�H��(�H�| ���  ������������H�AHÐ�������H�AH�H�D�Ð��H�H��H�Ð�����H9�t>H�L�IL�L�RI9�t,M9�L�YtOL�H�H�BH�AL�ZH�BL�AH�AL�B�M9�t8H�B�oABL�L�L�AH�AH�B��fD  �oRQH�L�	�H�y H�Bt(H��L�IL�Qt:      G�oJL�JL�RL�AIH�B�E1�H���{����oZYH�BH�AH�H�B    �  �L�JL�RH�AH�BH�H�A    �  ÐH�Ð�����������H�H�A    �  ÐVSH��(A�   H��H+H��H���C  H�H�H��([^Ð�����VSH��(H��H�	H��H)�HNI9�t%I)�H��H���  H�H�H��([^�f.�     H�^� H�H�H��([^Ð�����������VSH��(A�   H��H+H��H���  H�H�H��([^Ð�����VSH��(H��H�	H��H)�HNI9�t%I)�H��H���w  H�H�H��([^�f.�     H�^� H�H�H��([^Ð�����������SH�� L�IL9�H��w7I���tM��tI)�M9�MF��  H��H�� [�H�H�Q� H��H�� [�H�	y I��H�{y ��  ��H�Ð�����������VSH��(H��H��H���,���H��������H+KI��H9�rH��H��H��([^�  H��y ��  ���������H��(H��������H+AI9�w	H��(��  H�wy �T�  ����L�BH���  ����H��(L�RH�L��L)�L9�IG�M9�wL�I��H��(�  H�+y M��H�x �.�  ��������������H��(H��H�L�@H��������H+AI9�w	H��(�F  H��x ��  ����������H��8I��H�QE��D�D$ E1��t���H��8Ð��������������SH�� L�IH��H��H�H�L�CL9�tbL9�t=H�H�KH��L�HH�HH�KH�Ht4H�L�KH�C    � H�� [�f�     H�H�SH�PH�SH�PL�L����D  H��H��H�D$0�   ;      H�H�D$0묐�����VSH��8H��H��H���<���L�CI��1�H�D$ H���F���H��8[^Ð��������������H��8L�D$ L�AI��1�����H��8Ð���SH�� H���  H��H�� [Ð���������H��8L�RH�L��L)�L9�IG�M9�wN�H�D$ L�A1�����H��8�H�,w M��H�1v �D�  ����H��8H�BL�AH�D$ L�
1�����H��8�H��8E��I��1�D�D$ L�A����H��8�VSH��8A�   H��H+E��H��D�D$ E1�H������H�H�H��8[^Ð���������VSH��8H��H+E��H��D�L$ M��E1�H���J���H�H�H��8[^Ð������������H��8H+H�AM�M�@H9�wL�D$ E1������H��8�H�7u I��I��H��u �=�  �������������VSH��8A�   H��H+E��H��D�D$ E1�H������H�H�H��8[^Ð���������H��8H+E��D�L$ M��E1������H��8Ð��������������WVSH��0H��L��H��L������L�NL9�wH�D$ I��E1�H��H�������H��0[^_�H�$u I��H�Xt �k�  �����������H��8H�AH9�wL�L$ M��E1�����H��8�H�t I��I��H��t �%�  �����H��8H�AM�PM�H9�wL�T$ E1��_���H��8�H��s I��I��H��t ���  �H��(M�XM��L�L$PL��L)�L9�IG�M9�M�wL�AM�L9�w*E1�H�D$PH��(�����H�,t M��M��H�rs ��  H�fs M��I��H�t �l�  ������������H��8H�AH9�E��wD�L$ M��E1������H��8�H�s I��I��H��s<       �!�  �H��8H+H�AM)�H9�wL�L$ M��E1��]����H��8�H�h} I��I��H�C} ���  ��������������L�BLH��L�Ð�E1��   ��������H��8H�AH9�rvH�H�Q� H��8ÐH)�E��D�D$ I��E1�H���&����H��8�H�Ð�����������I��tM��u�@ �������Ð����I��tM��u�@ �Ӑ����Ð����H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�D���H��r M��I��H��q ���  �����������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�����H�'r M��I��H�Xq �k�  �����������H��8L�QM�YM�	H��H+I)�L��H)�I9�LG�L9�wL�\$ H������H��8�H��q M��I��H��p ��  �����������UWVSH��8H��L��H��L��L���$���L�NH��H)�H+I��L��H)�H9�LG�L9�wH��H�D$ I��H������H��8[^_]�H�Iq I��H�}p ��  ����������������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(����H��p M��I��H�p �+�  �����������H��(L�QH��H+I)�L��H)�I9�LG�L9�wH��H��(�Q���H��p M��I��H��o ���  ��������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�����H�7p M��I��H�ho �{�  �����������H��8L�QM�M�IH��H+I)�L��H)�I9�LG�L9�wL�L$ H��M������H��8�H=      ��o M��I��H�o ��  ��������D�T$(H��H+D�T$(I)������������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(����H�y M��I��H�y ��  �����������UWVSH��8H��L��H��L��L��贌��L�NH��H)�H+I��L��H)�H9�LG�L9�wH��H�D$ I��H������H��8[^_]�H��x I��H��x � �  ����������������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�4���H�-x M��I��H�8x ��  �����������H��(L�QH��H+I)�L��H)�I9�LG�L9�wH��H��(�����H��w M��I��H��w �h�  ��������H��8L�QM�YM�	H��H+I)�L��H)�I9�LG�L9�wL�\$ H������H��8�H�}w M��I��H��w ��  �����������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�$���H�w M��I��H�(w ��  �����������H��(L�YL�T$PH��H+I)�L��M)�H)�I9�LG�L9�wH��L�T$PH��(�����H��v M��I��H��v �K�  �����������D�T$(H��H+D�T$(I)�������������UWVSH��8H��L��L��H��L���D���L�OL��H)�H9�HF�L9�I��wH�D$ I��H��H���8���H��8[^_]�H�rl I��H��k ��  ���������H��(L�QL��H)�L9�LF�L9�w	H��(�����H�nk I��M��H�#l �t�  ����H��8L�QM�YM�	L��H)�L9�LF�L9�wL�\$ ����H��8�H�!k I>      ��M��H��k �'�  �������VSH��(I�YL�\$`H�t$hM�	H��L)�H9�HG�I9�w)M�L�YM��I)�M9�MF�L9�w)H�D$`H��([^�.���H�qk I��M��H��j ��  H��j I��M��H�Kk ��  ������������H��(L�QD�\$PL��H)�L9�LF�L9�wD�\$PH��(����H�Cj I��M��H��j �I�  ���������UWVSH��(H��H�IH�T$XH9�sH�L$XH��H�;H�sH9���   L�CI9�t9H��w@I9�r;H9�t)L�AI����   M��tH��H��興��H��� H�3H��([^_]�@ H�T$XH���C  H�;H��H�CL�@I��tOM��u*H9�tH���� H�D$XH�+H�CH��([^_]��     H��H�������� A�   �J���D  ��E ��     ��C�]��������VSH��(H�AN�L��I��M)�H��H�	t H��tI�H�I��t!L��蠇��H�H�CH)�H�C� H��([^�A��H�H�C��A�   H�AH�P������������������VSH��8H�AJ�4 H��H�	L�SL9�tSL�SL9�w*M��tH�I��tL�'���H�H��H�s�1 H��8[^�f�L�D$ I��H��E1�H���Z  H���D  A�   ��     ��H�벐�����ATUWVSH��0H9�H��H��t>H�9L�aH�rI9�tpL�AI9�r2H��tH��H�U tcH��I��舆��H�;H�s�7 H��0[^_]A\�f�H�T$(H��H�t$(�>   H�H��I9�t�� H�D$(H��H�;H�Ct��A�   � ��H�;롐�����H��(H�
H��xTL9�vM�L9�sM��x"I�HL�H��(�� f�?      H��H��(�  H��������H�       �H�H��(� H��f ���  ����H�QÐ����������AWAVAUATUWVSH��8H��$�   H��H�QL)�H��N�4M��L�iI��H�M)�L;)H�D$(��   L�AH�T$(H���(���H��H�;H��tH����   I��H��H���%���M��t/H��$�    t$H��$�   H�L5 ��   L��$�   L������M��t H�$�   J�7H��H�I��t4M���̄��I9�tH���O H�D$(H�+H�CH��8[^_]A\A]A^A_�f�����f�     ��E �`���D  A�   � ���D  A���t��������H��tH��u�@ A��I�Љ��2���f�D�Ð�����������UWVSH��8H�H�q��H��H�QH�~H9�tAH�QH9�w@�,0H�H�{�D0 H��8[^_]�H�D$    E1�E1�H��H���3���H��Ⱥ   뼐������H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�H�B    �B �f.�     �oBA�Ӑ����H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�H�B    �B �f.�     �oBAH�BH�AH�H�B    �  �VSH��(I������H�AH��H��H��H�tH���y���L�E1�H��H��H��([^�a����E1�H�AI�H��N�����������������H�AH�A    H��A Ð�����������E1�H�AH�H�L�BH��I����������E1�H�AH�H�L�BH��I���������H��(H�AH�H�BL�I9�wK�E1�M�H��(����H��d I��H�Lc �_�  ���������������H��(H�A@      H�H�BL�I9�wK�L)�L9�IG�E1�L�H��(�[���H�nd I��H��b ��  �����H��(H�AH�H�BL�I9�wK�L)�L9�IG�E1�L�H��(����H�9d I��H��b ��  �����E1�H�L�AL�L�BH��I����������H�AH�A    H��A Ð�����������H�AE��H������E1�H�AH�������E1�H�AH������E1�H�AH��1����H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�H�B    �B �f.�     �oBA�Ӑ����H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�H�B    �B �f.�     �oBAH�BH�AH�H�B    �  �VSH��(I������H�AH��H��H��H�tH�����L�E1�H��H��H��([^�����E1�H�AI�H��n�����������������H�AH�A    H��A Ð�����������E1�H�AH�H�L�BH��I����������E1�H�AH�H�L�BH��I����������H��(H�AH�H�BL�I9�wK�E1�M�H��(�����H��a I��H�l` ��  ���������������H��(H�AH�H�BL�I9�wK�L)�L9�IG�E1�L�H��(�{���H��a I��H�` �%�  �����H��(H�AH�H�BL�I9�wK�L)�L9�IG�E1�L�H��(�+���H�Ya I��H��_ ���  �����E1�H�L�AL�L�BH��I����������H�AH�A    H��A Ð�����������H�AE��H������E1�H�AH������E1�H�AH������E1�H�AH��Q����A      H�H�AH9�tH���| Ð����������H�H�AH9�tH���\ Ð����������SH�� L�IH��H��H�H�L�CI9�tbI9�t=H�H�KH��L�HH�HH�KH�Ht4H�L�KH�C    � H�� [�f�     H�H�SH�PH�SH�PL�L����D  H��H��H�D$0�`���H�H�D$0묐�����VSH��8H��H��H���|��L�CI��1�H�D$ H������H��8[^Ð��������������SH�� H������H��H�� [Ð���������SH��0H�BL�AH�D$ L�
H��1��Q���H��H��0[Ð�������SH��0A�   L�A��H�ˉT$ 1��p���H��H��0[Ð������H�H�Ð��������VSH��(H��H��H����{��H��������H+KI��H9�wH��H��H��([^����H�L^ �)�  ���������L�BH���������H��(H��H�L�@H��������H+AI9�w	H��(�f���H��] �ڼ  ����������UWVSH��8H�H�q��H��H�QH�~H9�tOH�QH9�w&@�,0H�H�{�D0 H��H��8[^_]�f.�     H�D$    E1�E1�H��H������H�뻐�   뮐��������H�	� ��������H�H�AH9�tH��� Ð����������AWAVAUATUWVSH��HH��������?H��$�   H��H�IL�L��H)�H9���  H�I��M)�L�CN�$)L9���  L�CM9��^  L�4PI��H�I)�@��H9���!�L9�vp@��t+I�~I��I�v�K  O�?L��$�   �Pz��L��$�   H��tH���  L�6L��L���2z��H�1�L�cfB�`H��H��H[^_]A\A]A^A_�H�HI9�wB      �H���  H9���   H����   L�6L��L��L��$�   M��L�T$8��y��@��L�T$8L��$�   t�f.�     I�~I��K���   O�?L��$�   �y��L��$�   H9��J���H�,6I�~I�)H9���   L9���   K�iH���  I��L���Ey������H�t$ I��H���  �����A�fA�������f������ A�   �^���D  A�fA�@���j���L�6�6���fD  H��t�I��L��L����x�������    �f��0���D  H��L)�I��I��I��t;M��tI��L��L���x��I�.L)�I�>H��t!H���?���L�6�hx���1���A�fA����f������fA�����H��] �V�  ����������H)�H������@H��   �M�ÐH�QÐ����������H�Ð�����������H�Ð�����������H�Ð�����������H�Ð�����������WVSH�� H��H��H�T$HD��D��w5H�H��t1�H��tED  f�HH��H9�u�1�H�Vf�PH�� [^_ÐH�T$HE1���  H�T$HH�H�V�D  f�8�Ȑ����������WVSH��0L��H��H��H)�H��H��H��H�T$(w,H��H�u�f�1�H�Vf�PH��0[^_�H��t��@ H�T$(E1��C  H�T$(H�H�VH��I��H����v��H�T$(H�벐��������������WVSH��0L��H��H��H)�H��H��H��H�T$(w,H��H�u�f�1�H�Vf�PH��0[^_�H��t��@ H�T$(E1��  H�T$(H�H�VH��I��H���9v��H�T$(H�벐��������������WVSH��0H��H��H��C      uM��u}L��H)�H��H��H��H�T$(w2H��H�u�f�1�H�Vf�PH��0[^_ÐH��t��%f�     H�T$(E1�H���  H�T$(H�H�VH��I��H���u��H�T$(H��H��[ 萵  ����������������WVSH��0H��H��H��uM��u}L��H)�H��H��H��H�T$(w2H��H�u�f�1�H�Vf�PH��0[^_ÐH��t��%f�     H�T$(E1�H���`  H�T$(H�H�VH��I��H����t��H�T$(H��H��Z ��  ����������������H�AÐ����������H�H�Q1�f�PÐ�I)�L��H��H��tH��u��t��fD  �f�Ð��������I)�L��H��H��tH��u��Vt��fD  �f�Ð��������I)�L��H��H��tH��u��&t��fD  �f�Ð��������I)�L��H��H��tH��u���s��fD  �f�Ð��������H��(H�AH9t#H�AH9Ar	H��(�@ 1��)  �H��(� �   ��H���q �H��(� �������AUATUWVSH��8H��������?D��$�   I��H�QL�H��L��D��H)�I9���   H�AL��L�	L)�H�I9���   H�AH9�rqK�(H)�t*I9�t%K�iH��N�@H�X��   L�L����r��L�H��tK�i1�H��t]f�,BH��H9�u�1�H�~fA�yH��H��8[^_]A\A]�D  E1�H�\$ L��H���  H��L�t�� �   �`���fD  fD�"�f.�     A�H��f�t��v���H��W 胳  ���H��Ð�����������E�������������H��(L�AL9�sH�H�PH��(�H�W �k�  ���D      ��������H�QH�H�PÐ���H�QH�H�DP�Ð��H�H��H�Ð�����H9�t>H�L�IL�L�RI9�t,M9�L�YtOL�H�H�BH�AH�BL�ZL�AH�AL�B�M9�H�Bt4L�J�oABL�L�AL�L�I��fD  �oRQH�L�	�H�y t(H��L�IL�QtK�oJL�JL�RL�AIH�B�E1�H��t��oZYH�BH�AH�1�H�B    f��fD  L�JL�RH�AH�BH�1�H�A    f�Ð��������������H�Ð�����������1�H�H�A    f�Ð��������������VSH��(A�   H��H+H��H��H���   H�H�H��([^Ð��VSH��(H��H�	H��H��L�KH)�J�IH��H��I9�tI)�H��I���  H�H�H��([^�H�S1�f�H��([^Ð������������VSH��(A�   H��H+H��H��H���p  H�H�H��([^Ð��VSH��(H��H�	H��H��L�KH)�J�IH��H��I9�tI)�H��I���*  H�H�H��([^�H�S1�f�H��([^Ð������������SH�� L�IL9�H��w9I���tM��tI)�M9�MF���  H��H�� [�H�H�Q1�f�PH��H�� [�H��S I��H�YT �p�  ����������������H�Ð�����������VSH��(H��H��H���$n��H��������?H+KI��H9�wH��H��H��([^��  H�|T �ٯ  ���������H��(H��������?H+AI9�w	H��(�  H�GT 褯  ����L�BH��  ����H��(L�RH�L��L)�L9�IG�M9�wJ�BI��H��(�S  H��S M��H��R �}�  �������������E      H��(H��H�L�@H��������?H+AI9�w	H��(�  H��S �
�  ����������H��8I��H�QE��D�D$ E1��4���H��8Ð��������������SH�� L�IH��H��H�H�L�CL9�tUL9�L�[L�St5H��L�HH�L�XL�Pt,H�L�K1�H�C    f�
H�� [��    H�L�XL�PL�L����H��H��H�D$0��  H�H�D$0빐��VSH��8H��H��H���Dl��L�CI��1�H�D$ H�������H��8[^Ð��������������H��8L�D$ L�AI��1������H��8Ð���SH�� H���S  H��H�� [Ð���������H��8L�RH�L��L)�L9�IG�M9�wN�BH�D$ L�A1��o���H��8�H�R M��H�Q 褳  ����H��8H�BL�AH�D$ L�
1��5���H��8�H��8E��I��1�D�D$ L�A����H��8�VSH��8A�   H��H+E��H��D�D$ E1�H��H���T���H�H�H��8[^Ð������VSH��8H��H+E��H��D�L$ M��E1�H��H������H�H�H��8[^Ð���������H��8H+H�AM�M�@H��H9�wL�D$ E1��i����H��8�H�P I��I��H��P 蚲  ����������VSH��8A�   H��H+E��H��D�D$ E1�H��H������H�H�H��8[^Ð������H��8H+E��H��D�L$ M��E1��R����H��8Ð�����������WVSH��0H��L��H��L����i��L�NL9�wH�D$ I��E1�H��H������H��0[^_�H�P I��H�8O �˱  �����������H��8H�AH9�wL�L$ M��E1��S���H��8�H��N I��I��H��O 腱  �����H��8H�AF      M�PM�H9�wL�T$ E1�����H��8�H��N I��I��H�pO �A�  �H��(L�\$PM��M�HM� L��L)�L9�IG�M9�wO�PL�AL9�w'E1�H�D$PH��(����H�O M��H�TN ��  H�HN M��I��H��N �ΰ  ��������������H��8H�AH9�E��wD�L$ M��E1�����H��8�H��M I��I��H��N 聰  �H��8H+H�AM)�H��I��H9�wL�L$ M��E1������H��8�H��T I��I��H��T �8�  ��������H��H�JH�H�JH�Ð�������������E1��   ��������H��8H�AH9�rvH�H�Q1�f�PH��8�H)�E��D�D$ I��E1�H��������H��8Ð��������������H�Ð�����������I��tM��u�@ M��8h���     �f�Ð��������I��tM��u�@ M�� h���     �f�Ð��������H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(����H�M M��I��H�LL �߮  ���������������H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(�8���H��L M��I��H��K �o�  ���������������H��8L�QM�YM�	H��H+I)�L��I��H��H)�I9�LG�L9�wL�\$ H�������H��8�H�AL M��I��H�rK ��  �����UWVSH��8H��H��L��L��L����e��L�NH��H)�H+I��I��L��H��H)�I9�LG�L9�wH��H�D$ I��H���Y���H��8[^_]�H��K I��H��J 芭  ����������G      H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(�����H�[K M��I��H��J ��  ���������������H��(L�QH��H+I)�L��I��H��H)�I9�LG�L9�wH��H��(����H��J M��I��H�/J �¬  ��H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(�(���H��J M��I��H��I �_�  ���������������H��8L�QM�M�IH��H+I)�L��I��H��H)�I9�LG�L9�wL�L$ H��M�������H��8�H�.J M��I��H�_I ��  ���D$(I)�H+�D$(I��H�������������H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(�8���H��O M��I��H��O �o�  ���������������UWVSH��8H��H��L��L��L���,c��L�NH��H)�H+I��I��L��H��H)�I9�LG�L9�wH��H�D$ I��H������H��8[^_]�H�YO I��H�gO ��  ����������H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(�H���H��N M��I��H��N ��  ���������������H��(L�QH��H+I)�L��I��H��H)�I9�LG�L9�wH��H��(�����H��N M��I��H��N �"�  ��H��8L�QM�YM�	H��H+I)�L��I��H��H)�I9�LG�L9�wL�\$ H������H��8�H�7N M��I��H�BN �ũ  �����H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wHH      ��L�T$PH��(�(���H��M M��I��H��M �_�  ���������������H��(H�D$PL�YL)�I)�H��I��I��H��H+L��H��H)�I9�LG�L9�wH��L�T$PH��(����H�aM M��I��H�lM ��  ����������������D$(I)�H+�D$(I��H�������������UWVSH��8H��L��L��H��L���`��L�OL��H)�H9�HF�L9�I��wH�D$ I��H��H���(���H��8[^_]�H��F I��H��E �Y�  ���������H��(L�QL��H)�L9�LF�L9�w	H��(�����H��E I��M��H�CF ��  ����H��8L�QM�YM�	L��H)�L9�LF�L9�wL�\$ ����H��8�H�AE I��M��H��E �ǧ  �������VSH��(I�YL�\$`H�t$hM�	H��L)�H9�HG�I9�w*O�YL�YM��I)�M9�MF�L9�w)H�D$`H��([^����H��E I��M��H��D �T�  H��D I��M��H�jE �;�  �����������H��(L�QD�\$PL��H)�L9�LF�L9�wD�\$PH��(�"���H�cD I��M��H�E ��  ���������UWVSH��(H��H�IH�T$XH9�sH�L$XH��H�;H�sH9���   L�CI9�t=H��w@I9�r;H9�t-H��H����   H��tL�	H��H���$_��H����  H�3H��([^_]�H�T$XH���c  H�;H��H�CL�@I��tOM��u*H9�tH���m�  H�D$XH�+H�CH��([^_]��     M�H��H���^����A�   �J���D  �f�E ��    �f�C�`�������VSH��(H�AH��L��J�I��L�I)�t%H��t M�II��I�Qt.M�L���;^��L�I      H�CH)�1�H�CfA�AH��([^��    A�f��ې������A�   H�AH�P��}����������������VSH��8H��H�IH�L�SJ�4L9�tSL�SL9�w.M��tH�HI��tKM��]��H�1�H�sf�pH��H��8[^�L�D$ I��E1�H��H���f  H��ѐA�   ��     �f�븐�������ATUWVSH��0H9�H��H��tAH�9L�aH�rI9�t{L�AI9�r3L�6H��tH��H�U toH���]��H�;1�H�sf�wH��0[^_]A\�H�T$(H��H�t$(�M   H�H��I9�t�m�  H�D$(H�;L�6H��H�Ct��fD  A�   ��     �f�딐�������H��(H��������?H�H9�w>L9�v+M�L9�s#I9�vH�
H�       �H��(�2�  f�L�L��H�L H��(��  H��@ �`�  ����������������H�QÐ����������AWAVAUATUWVSH��8H��$�   H��H�QL)�H��N�4M��L�aI��H�M)�L;!H�D$(��   L�AH�T$(H���(���H��H�;H��tH����   L�6H��H���[��M��t3H��$�    t(H��$�   H�Lu ��   H��$�   L��L� �l[��M��t!H�$�   J�wI��H�Lu t4O�D- �F[��I9�tH�����  H�D$(H�+H�CH��8[^_]A\A]A^A_��f���@ �f�E �`���@ A�   � ���D  A�f��x�������H��E��tH��t1�fD�AH��H9�u�ÐfD�Ð����������UWVSH��8H�H�q��H��H�QH�~H9�t@H�QH9�w1�f�,pH�{f�TpH��8[^_]�H�D$    E1�E1�H��H���4���H��ɺ   �J      ��������H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�1�H�B    f�B��     �oBA�Ӑ����H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�1�H�B    f�B��     �oBAH�BH�AH�H�B    1�f�Ð�������������SH��0I������H�AH��H��H�tH��H�T$(�X��H�T$(L�BE1�H��H��0[�������������������E1�H�AN�BH�������������������H�AH�A    H�1�f�AÐ���������E1�H�AH�H�H�RL�PH���c������E1�H�AH�H�H�RL�PH���s������H��(L�JH�AM9�H�H�wJ�@L��E1�L)�L�BH��(�_���H��> H�)= 輟  ������������H��(H�AH�H�BL�I9�wK�BL)�L9�IG�E1�L�BH��(����H�N> I��H��< �e�  �����H��(H�AH�H�BL�I9�wK�BL)�L9�IG�E1�L�BH��(����H�> I��H��< ��  �����E1�H�H�RL�AL�L�PH���������H�AH�A    H�1�f�AÐ���������H�AE��H�����E1�H�AH������E1�H�AH��1����E1�H�AH�������H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�1�H�B    f�B��     �oBA�Ӑ����H�AH�L�H�BL9�t-L�L�BL�AL�BL�AH�1�H�B    f�B��     �oBAH�BH�AH�H�B    1�f�Ð�������������SH��0I������H�AH��H��H�tH��H�T$(�U��H�T$(L�K      BE1�H��H��0[�������������������E1�H�AN�BH�������������������H�AH�A    H�1�f�AÐ���������E1�H�AH�H�H�RL�PH���c������E1�H�AH�H�H�RL�PH���s������H��(L�JH�AM9�H�H�wJ�@L��E1�L)�L�BH��(�_���H��; H�): 輜  ������������H��(H�AH�H�BL�I9�wK�BL)�L9�IG�E1�L�BH��(����H�N; I��H��9 �e�  �����H��(H�AH�H�BL�I9�wK�BL)�L9�IG�E1�L�BH��(����H�; I��H��9 ��  �����E1�H�H�RL�AL�L�PH���������H�AH�A    H�1�f�AÐ���������H�AE��H�����E1�H�AH������E1�H�AH��1����E1�H�AH�������H�H�AH9�tH����  Ð����������H�H�AH9�tH����  Ð����������SH�� L�IH��H��H�H�L�CI9�tUI9�L�[L�St5H��L�HH�L�XL�Pt,H�L�K1�H�C    f�
H�� [��    H�L�XL�PL�L����H��H��H�D$0����H�H�D$0빐��VSH��8H��H��H���R��L�CI��1�H�D$ H���F���H��8[^Ð��������������SH�� H�������H��H�� [Ð���������SH��0H�BL�AH�D$ L�
H��1������H��H��0[Ð�������SH��0A�   L�A��H�ˉT$ 1��0���H��H��0[Ð������H�H�PÐ�������VSH��(H��H��H����Q��H��������?H+KI��H9�wH��H��H��([^�u���H�8 �y�  �L      ��������L�BH��T�������H��(H��H�L�@H��������?H+AI9�w	H��(�&���H��7 �*�  ����������UWVSH��8H�H�q��H��H�QH�~H9�tCH�QH9�w1�f�,pH�{f�TpH��H��8[^_]�H�D$    E1�E1�H��H������H��ƺ   뺐����ATUWVSH�� L�%_� 1�M��L�!H��H�����A�6���H�CH�� �   H��H�H�=N* ��� ��tH�=>* �   H����� ��uH�� [^_]A\�f�     H�sH���t���E1�H��H�������H�� [^_]A\�H��L�#H���L���H���t���H���̨��H��H���a���H��蹨�����������ATUWVSH�� L�%� 1�H�*M��L�!H�����A�V���H�CH�;� �   H��H�H�=n) ��� ��tH�=^) �   H����� ��uH�� [^_]A\�f�     H�sH��蔚��E1�H��H���&����H�� [^_]A\�H��L�#H���l���H��蔚��H������H��H��聚��H���٧�����������ATUWVSH�� L�%�� 1�M��L�!H��H�����A�v���H�CH�[� �   H��H�H�=�( ��� ��tH�=~( �   H����� ��uH�� [^_]A\�f�     H�sH��贙��E1�H��H���F����H�� [^_]A\�H��L�#H��茙��H��贙��H������H��H��衙��H����������������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A薘��H�CH�{� �   H��H�H�=�' ��� ��tH�=�' �   H����� ��uH�� [^_]A\�f�     H�sH���Ԙ��E1�HM      ��H���f����H�� [^_]A\�H��L�#H��謘��H���Ԙ��H���,���H��H�������H���������������SH�� H��� H�H��H�I�e���H��荘��H��H�� [�p�  SH�� H��� H�H��H�I�5���H��H�� [�X�����������SH�� H��� H�H��H�I����H��H�� [�(�����������ATUWVSH�� L�%�� 1�M��L�!H��H�����A�&���H�CH�K� �   H��H�H�=) ��� ��tH�=�( �   H����� ��uH�� [^_]A\�f�     H�sH���d���E1�H��H��������H�� [^_]A\�H��L�#H���<���H���d���H��輤��H��H���Q���H��詤�����������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A�F���H�CH�k� �   H��H�H�=.( ��� ��tH�=( �   H����� ��uH�� [^_]A\�f�     H�sH��脖��E1�H��H�������H�� [^_]A\�H��L�#H���\���H��脖��H���ܣ��H��H���q���H���ɣ�����������ATUWVSH�� L�%�� 1�M��L�!H��H�����A�f���H�CH��� �   H��H�H�=N' ��� ��tH�=>' �   H����� ��uH�� [^_]A\�f�     H�sH��褕��E1�H��H���6����H�� [^_]A\�H��L�#H���|���H��褕��H�������H��H��葕��H���������������ATUWVSH�� L�%�� 1�H�*M��L�!H�����A膔��H�CH��� �   H��H�H�=n& ��� ��tH�=^& �   H����� ��uH�� [^_]A\�fN      �     H�sH���Ĕ��E1�H��H���V����H�� [^_]A\�H��L�#H��蜔��H���Ĕ��H������H��H��豔��H���	������������SH�� H�� H�H��H�I�U���H���}���H��H�� [�`�  SH�� H��� H�H��H�I�%���H��H�� [�H�����������SH�� H��� H�H��H�I�����H��H�� [������������UWVSH��(H�=f" H��L��H����   H��� �   H��H���� ��tH�=6" �   H����� ��uH��([^_]� H�sH���t���E1�H��H�������H��([^_]�H��H��H�?� H��G���H���o���H���Ǡ���������H��H�����������UWVSH��(H�=�! H��L��H���   H��� �   H��H���� ��tH�=v! �   H����� ��uH��([^_]� H�sH��贒��E1�H��H���F����H��([^_]�H��H��H�� H�臒��H��诒��H�������������H�������������SH�� H�D� H�H��H�I�E���H���m���H��H�� [�P�  SH�� H�� H�H��H�I����H��H�� [�8�����������SH�� H��� H�H��H�I����H��H�� [������������UWVSH��(H�=&# H��L��H���   H��� �   H��H���� ��tH�=�" �   H����� ��uH��([^_]� H�sH���d���E1�H��H��������H��([^_]�H��H��H�o� H��7���H���_���H��跞���������H��H�����������UWVSH��(H�=f" H��L��H����  H��� �   H��H��O      ��� ��tH�=6" �   H����� ��uH��([^_]� H�sH��褐��E1�H��H���6����H��([^_]�H��H��H��� H��w���H��蟐��H��������������H�������������SH�� H�t� H�H��H�I�5���H���]���H��H�� [�@�  SH�� H�D� H�H��H�I����H��H�� [�(�����������SH�� H�� H�H��H�I�Տ��H��H�� [�������������UWVSH��81�M��H��H�A    H����1҉AH�� H��N  H��� �   H��H�H�=
 ��� ��tH�=� �   H����� ��uH��8[^_]��    H�t$(E1�H��H���͎��H�T$(H����  H�������H��8[^_]�H��H���"  H��苜��H��H��� ���H���x�����������UWVSH��81�H�*M��H�A    H����1҉AH�&� H��n  H��� �   H��H�H�=* ��� ��tH�= �   H����� ��uH��8[^_]��    H�t$(E1�H��H������H�T$(H���   H���8����H��8[^_]�H��H���#!  H��諛��H��H���@���H��蘛����������UWVSH��81�M��H��H�A    H����1҉AH�F� H��  H�� �   H��H�H�=J ��� ��tH�=: �   H����� ��uH��8[^_]��    H�t$(E1�H��H������H�T$(H���   H���X����H��8[^_]�H��H���C   H���˚��H��H���`���H��踚����������UWVSH��81�H�*M��H�A    H����1҉AH�f� H��  H�7�P       �   H��H�H�=j ��� ��tH�=Z �   H����� ��uH��8[^_]��    H�t$(E1�H��H���-���H�T$(H���@  H���x����H��8[^_]�H��H���c  H������H��H��而��H���ؙ����������SH�� H��� H��H��)  H��H�� [�<�  ������������H�Y� H��  �H�I� H���  �UWVSH��81�M��H��H�A    H����1҉AH��� H��  H�W� �   H��H�H�=
 ��� ��tH�=� �   H����� ��uH��8[^_]��    H�t$(E1�H��H�������H�T$(H���  H���H����H��8[^_]�H��H���!  H��軘��H��H���P���H��記����������UWVSH��81�H�*M��H�A    H����1҉AH��� H��.  H�w� �   H��H�H�=* ��� ��tH�= �   H����� ��uH��8[^_]��    H�t$(E1�H��H������H�T$(H����  H���h����H��8[^_]�H��H����   H���ۗ��H��H���p���H���ȗ����������UWVSH��81�M��H��H�A    H����1҉AH��� H��N  H��� �   H��H�H�=J ��� ��tH�=: �   H����� ��uH��8[^_]��    H�t$(E1�H��H���=���H�T$(H����  H��舉���H��8[^_]�H��H����  H�������H��H��萉��H��������������UWVSH��81�H�*M��H�A    H����1҉AH��� H��n  H��� �   H��H�H�=j ��� ��tH�=Z � Q        H����� ��uH��8[^_]��    H�t$(E1�H��H���]���H�T$(H���   H��計���H��8[^_]�H��H���  H������H��H��谈��H��������������SH�� H�� H��H���  H��H�� [�l�  ������������H��� H��  �H��� H��  �1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������1�M�����AH��� H�Ð���������SH�� H��� H��H�蹇��H��H�� [��  ������������H�y� H�鑇���H�i� H�遇���1�M�����AH��� H�Ð���������1�M�����AH�n� H�Ð���������1�M�����AH�N� H�Ð���������1�M�����AH�.� H�Ð���������SH�� H�4� H��H�����H��H�� [���  ������������H�	� H�������H��� H�鱆���UWVSH��81�M��H��H�A    H����E1�1҉AH��� H��;���H��� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H��荅��H�T$(E1�H���͈��H���Յ���H��8[^_]�H��H��� ���H���H���H��H���݅��H���5��������UWVSH��81�H�*M��H�A    H����E1�1҉AH�� H��[���H�� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H��譄��H�T$(E1�H������H����R      ����H��8[^_]�H��H���@���H���h���H��H�������H���U��������UWVSH��81�M��H��H�A    H����E1�1҉AH�#� H��{���H�4� �   H��H�H�= ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���̓��H�T$(E1�H������H�������H��8[^_]�H��H���`���H��舑��H��H������H���u��������UWVSH��81�H�*M��H�A    H����E1�1҉AH�C� H�蛆��H�T� �   H��H�H�=' ��� ��tH�= �   H����� ��uH��8[^_]�@ H�t$(E1�H��H������H�T$(E1�H���-���H���5����H��8[^_]�H��H��耉��H��訐��H��H���=���H��蕐�������SH�� H��� H��H��I���H��H�� [���  ������������H�y� H��!����H�i� H������UWVSH��81�M��H��H�A    H����E1�1҉AH��� H��+���H��� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H��轁��H�T$(E1�H��轈��H�������H��8[^_]�H��H������H���x���H��H������H���e��������UWVSH��81�H�*M��H�A    H����E1�1҉AH��� H��K���H��� �   H��H�H�= ��� ��tH�= �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���݀��H�T$(E1�H���݇��H���%����H��8[^_]�H��H���0���H��蘎��H��H���-S      ���H��腎�������UWVSH��81�M��H��H�A    H����E1�1҉AH��� H��k���H��� �   H��H�H�=7 ��� ��tH�=' �   H����� ��uH��8[^_]�@ H�t$(E1�H��H������H�T$(E1�H�������H���E����H��8[^_]�H��H���P���H��踍��H��H���M���H��襍�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�� H�苆��H��� �   H��H�H�=W ��� ��tH�=G �   H����� ��uH��8[^_]�@ H�t$(E1�H��H�����H�T$(E1�H������H���e���H��8[^_]�H��H���p���H���،��H��H���m��H���Ō�������SH�� H�D� H��H��9���H��H�� [�,�  ������������H�� H������H�	� H������UWVSH��81�M��H��H�A    H����E1�1҉AH�#� H�����H�4� �   H��H�H�=� ��� ��tH�=� �   H����� ��uH��8[^_]�@ H�t$(E1�H��H����}��H�T$(E1�H��譈��H���5~���H��8[^_]�H��H������H��訋��H��H���=~��H��蕋�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�C� H��;���H�T� �   H��H�H�= ��� ��tH�= �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���}��H�T$(E1�H���͇��H���U}���H��8[^_]�H��H���0���H���Ȋ��H��H���]}��H��赊�������UWVSH��81�M��H��H�A    T      H����E1�1҉AH�c� H��[���H�t� �   H��H�H�=7 ��� ��tH�=' �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���-|��H�T$(E1�H������H���u|���H��8[^_]�H��H���P���H������H��H���}|��H���Չ�������UWVSH��81�H�*M��H�A    H����E1�1҉AH��� H��{���H��� �   H��H�H�=W ��� ��tH�=G �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���M{��H�T$(E1�H������H���{���H��8[^_]�H��H���p���H������H��H���{��H������������SH�� H�� H��H��9���H��H�� [�\�  ������������H��� H������H��� H������UWVSH��81�M��H��H�A    H����E1�1҉AH�û H�����H�Կ �   H��H�H�=' ��� ��tH�= �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���z��H�T$(E1�H��譈��H���ez���H��8[^_]�H��H������H���؇��H��H���mz��H���Ň�������UWVSH��81�H�*M��H�A    H����E1�1҉AH�� H��;���H��� �   H��H�H�=G ��� ��tH�=7 �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���=y��H�T$(E1�H���͇��H���y���H��8[^_]�H��H���0���H�������H��H���y��H�����������UWVSH��81�M��H��H�A    H����E1�1҉AH�� H��[���H�� �  U       H��H�H�=g
 ��� ��tH�=W
 �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���]x��H�T$(E1�H������H���x���H��8[^_]�H��H���P���H������H��H���x��H�����������UWVSH��81�H�*M��H�A    H����E1�1҉AH�#� H��{���H�4� �   H��H�H�=�	 ��� ��tH�=w	 �   H����� ��uH��8[^_]�@ H�t$(E1�H��H���}w��H�T$(E1�H������H����w���H��8[^_]�H��H���p���H���8���H��H����w��H���%��������SH�� H��� H��H��9���H��H�� [錽  ������������H�Y� H������H�I� H������SH�� 1�M��H��H�T$8���AH��� H�H�L$8�v��H�CH�� [Ð���������VSH��(1�H��H�����AH�U� H��=v��H�CH��([^�H��H����v��H���O������������������SH�� 1�M��H��H�T$8���AH�� H�H�L$8�v��H�CH�� [Ð���������VSH��(1�H��H�����AH�Ż H��u��H�CH��([^�H��H���gv��H��迃�����������������SH�� H��� H�H��H�I�v��H���-v��H��H�� [��  SH�� H�T� H�H��H�I��u��H��H�� [��u����������SH�� H�$� H�H��H�I�u��H��H�� [��u����������SH�� 1�M��H��H�T$8���AH�!� H�H�L$8��t��H�CH�� [Ð���������VSH��(1�H��H�����AH�� H��t��H�CH��([^�H��H���Gu�V      �H��蟂�����������������SH�� 1�M��H��H�T$8���AH��� H�H�L$8�dt��H�CH�� [Ð���������VSH��(1�H��H�����AH�U� H���s��H�CH��([^�H��H���t��H���������������������SH�� H�� H�H��H�I�Ut��H���}t��H��H�� [�`�  SH�� H�� H�H��H�I�%t��H��H�� [�Ht����������SH�� H��� H�H��H�I��s��H��H�� [�t����������VSH��(1�M��H�����AH��� H��s��H�CH��([^�H��H����s��H���/������������������VSH��(1�H��H�����AH�e� H���r��H�CH��([^�H��H���s��H���߀�����������������VSH��(1�M��H�����AH�� H��}r��H�CH��([^�H��H���7s��H��菀�����������������VSH��(1�H��H�����AH�Ÿ H��-r��H�CH��([^�H��H����r��H���?������������������SH�� H��� H�H��H�I�r��H���r��H��H�� [鐸  SH�� H�T� H�H��H�I�Ur��H��H�� [�xr����������SH�� H�$� H�H��H�I�%r��H��H�� [�Hr����������VSH��(1�M��H�����AH�%� H��Mq��H�CH��([^�H��H���r��H���_�����������������VSH��(1�H��H�����AH�շ H���p��H�CH��([^�H��H���q��H��������������������VSH��(1�M��H�����AH��� H��p��H�CH��([^�H��H���gq��H���~�����������������W      VSH��(1�H��H�����AH�5� H��]p��H�CH��([^�H��H���q��H���o~�����������������SH�� H��� H�H��H�I�p��H����p��H��H�� [���  SH�� H�Ķ H�H��H�I�p��H��H�� [�p����������SH�� H��� H�H��H�I�Up��H��H�� [�xp����������SH�� H�AH��H����   H���  H�PH�CH�@    H�C�@  H�C�@H.H�C�@I,H�UA L� 1�A� H�S�LJH��H��$u�H�"A L� 1�A� H�S�LnH��H��u�H�CH�|�  H�z�  H�H(H�CH�@0   H�CH�P8H�CH�@@   H�� [ù�   �е  H��H �@    H�@    H�@    H�Q�@  H�1�H�@(    H�@0    H�@8    H�@@    f�PHƀ�    H�C������VSH��(1�M��H�QH����1҉AH�_� H������H��([^�H��H���o��H���\|��������������VSH��(1�M��H�A    H�����AH�� H��U����H��([^�H��H���n��H���
|������������VSH��(1�H��H�A    H����1҉AH��� H������H��([^�H��H���`n��H���{����������VSH��(1�M��H�QH����1҉AH�o� H������H��([^�H��H���n��H���l{��������������VSH��(1�M��H�A    H�����AH�� H��e����H��([^�H��H����m��H���{������������VSH��(1�H��H�A    H����1҉AH�˳ H������H��([^�H��H���pm��H����z����������VSH��(H�X      ��"   H��H��([^�4�  H��H���)�  H���z���VSH��(H��C H��H��H�H�IH��tH��PH��H��([^��l��H��H����l��H���Iz�����������SH�� H�AH��H����   H��= H�]�  �@  H�XH�@    �@H. , L�1ҐfA�f�LPLH��H��$u�H��= L�1�fA�f��P�   H��H��u�H��  H�@0   H�X(H��  H�X8H�@@   H�� [ù�   �a�  H�*E �@    H�@    H�@    H�Q�@  H�H�@(    H�@0    H�@8    H�@@    �@H    ƀ�    H�C�����VSH��(1�M��H�QH����1҉AH�?� H�������H��([^�H��H���k��H����x��������������VSH��(1�M��H�A    H�����AH�� H��u����H��([^�H��H���Bk��H���x������������VSH��(1�H��H�A    H����1҉AH��� H��#����H��([^�H��H����j��H���Hx����������VSH��(1�M��H�QH����1҉AH�O� H�������H��([^�H��H���j��H����w��������������VSH��(1�M��H�A    H�����AH��� H������H��([^�H��H���Rj��H���w������������VSH��(1�H��H�A    H����1҉AH��� H��3����H��([^�H��H��� j��H���Xw����������VSH��(H���"   H��H��([^�į  H��H��蹯  H���!w���VSH��(H��@ H��H��H�H�IH��tH��PH��H��([^�i��H��H���i��H����v�����������1�H�����AH�>�Y       H�Ð���������1�H�����AH�� H�Ð���������SH�� H�� H��H��i��H��H�� [���  ������������H�ٯ H���h���H�ɯ H���h���1�H�����AH�� H�Ð���������1�H�����AH�� H�Ð���������SH�� H�ԯ H��H��h��H��H�� [�l�  ������������H��� H��ah���H��� H��Qh���1�H�����AH�ޯ H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H���g��H��H�� [�ܭ  ������������H�y� H���g���H�i� H���g���1�H�����AH�~� H�Ð���������1�H�����AH�^� H�Ð���������SH�� H�D� H��H��ig��H��H�� [�L�  ������������H�� H��Ag���H�	� H��1g���1�H�����AH�� H�Ð���������1�H�����AH��� H�Ð���������SH�� H�� H��H���f��H��H�� [鼬  ������������H��� H��f���H��� H��f���1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H��If��H��H�� [�,�  ������������H�Y� H��!f���H�I� H��f���SH�� H��� H��H���e��H��H�� [�ܫ  ������������H�Y� H���e���SH�� H��� H��H��e��H��H�� [霫  ������������H�y� H��e���SH�� 1�M��H��H�T$8���AH�1� H�H�L$8�Z      �d��H�CH�� [Ð���������VSH��(1�H��H�����AH��� H��]d��H�CH��([^�H��H��> H��H�PH��	e��H���ar���VSH��(H���"   H��H��([^�Ԫ  H��H���ɪ  H���1r���VSH��(H��� H��H�H�I�d��H�M> H��H��H�H��([^�d��H��H�.> H��H�PH��d��H����q���������SH�� 1�M��H��H�T$8���AH�q� H�H�L$8�c��H�CH�� [Ð���������VSH��(1�H��H�����AH�5� H��=c��H�CH��([^�H��H��= H��H�PH���c��H���Aq���VSH��(H���"   H��H��([^鴩  H��H��詩  H���q���VSH��(H��� H��H�H�I�dc��H�== H��H��H�H��([^�xc��H��H�= H��H�PH��_c��H���p���������SH�� 1�M��H��H�T$8���AH��� H�H�L$8�b��H�CH�� [Ð���������VSH��(1�H��H�����AH�u� H��b��H�CH��([^�H��H����b��H���/p�����������������SH�� 1�M��H��H�T$8���AH�!� H�H�L$8��a��H�CH�� [Ð���������VSH��(1�H��H�����AH��� H��a��H�CH��([^�H��H���Gb��H���o�����������������SH�� H��� H�H��H�I��a��H���b��H��H�� [��  SH�� H�t� H�H��H�I�a��H��H�� [��a����������SH�� H�D� H�H��H�I�a��H��H�� [�a����������SH�� 1�M��H��H�T$8���AH�A� H�H�L$8��`��H�C[      H�� [Ð���������VSH��(1�H��H�����AH�� H��m`��H�CH��([^�H��H���'a��H���n�����������������SH�� 1�M��H��H�T$8���AH��� H�H�L$8�D`��H�CH�� [Ð���������VSH��(1�H��H�����AH�u� H���_��H�CH��([^�H��H���`��H����m�����������������SH�� H�4� H�H��H�I�5`��H���]`��H��H�� [�@�  SH�� H�� H�H��H�I�`��H��H�� [�(`����������SH�� H��� H�H��H�I��_��H��H�� [��_����������1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H��_��H��H�� [�|�  ������������H�y� H��q_���H�i� H��a_���1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H��	_��H��H�� [��  ������������H�i� H���^���H�Y� H���^���1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H��y^��H��H�� [�\�  ������������H�Y� H��Q^���H�I� H��A^���1�H�����AH��� H�Ð���������1�H�����AH�n� H�Ð���������SH�� H�T� H��H���]��H��H�� [�̣  ������������H�)� H���]���H�� H��]���SH�� H�d� H��H��9:  �   H��H�� [釣  �������H�9� H\      ��:  �ATUWVSH��0H�i@Hc�H�˃�~:�����u_�A ���A�A �E  E���  H�C0    H�C0H��0[^_]A\�A�   H��H���   H�D5 D���   H��0[^_]A\�D  D�fH�%3 D�D$(Ic�H��H����  D�D$(H����   H�O�H��H��H�    H���B�    H���u䋓�   ��~6D�J�1�I��I���     H���   L�L��L�LH��I9�u�H���   H��tTH9�tOH�D$(�%�  H�D$(H���!����     �C8    �����@ �C ���C�C �����H�g�  �O  f�H�������H���  ��N  ������������WVSH��0H�5�0 ���t��u
��H��0[^_�H�|$/H���/  H�H4 � H�, H�pH�1H��8�]��H��+ H�1H��8�]��H��+ H�1H��8�]��H�4 H�
, H�pH�1H��8�z]��H��+ H�1H��8�g]��H��+ H�1H��8�T]���   H�5H�  ��H��+ A�   A�   H����o��1���H��+ A�   A�   H���o���   ��H��+ A�   A�   H���o��H��0 H��+ H���3)  H�L0 H�U+ H���)  H�E0 H�N+ H���)  H�>0 H�7+ H����(  �   ��H�`+ A�   A�   H���s��1���H�!+ A�   A�   H����r���   ��H�+ A�   A�   H����r��H�$0 H��* H���1  H��/ H��* H���}1  H��/ H��* H���f1  H��/ H��* H���O1  H����  ��H��0[^_�H��H����  H�]      ���f������������WVSH�� H�Y(H��H�Ή�tD�CH����SH�H��u�H�� [^_�H���g�  肣  ��H��H��t�f����  �������������WVSH�� H�˹   H��D���&�  H�S(H�x�p�@    H�H�C(H�� [^_Ð����VSH��(H��H�I(H��u�H�褞  H��H��t�������A��t�H�F(    H��([^Ð��������������AVAUATUWVSH�� H�5+- �   ����tH�� [^_]A\A]A^�H�- �   L�%l�  � A��H��( H��H��0 H�K8H�C    L�hH�C    L�+H�C    H�C     H�C(    H�C0    �UY��H�.. H�{@1��CH����H�hH�+A��H�= ( I��H�O8L�/H�G    H�G    H�G    H�G     H�G(    H�G0    ��X��L�w@�   H�/�GH����A��H�=�' I��H�O8L�/H�G    H�G    H�G    H�G     H�G(    H�G0    �X��L�w@H�/�GH����H�=�, H�O�7  H�O1�H��L�5W. f���   HǇ�       HǇ�       HǇ�       HǇ       I�FH�I�F@HǇ      H�G�u"  H�-N, H�M��  1�Hǅ�       f���   H�MH��- Hǅ�       Hǅ       Hǅ      H�PH��@Hǅ      H�U H��& H�EH�E    ��!  H��+ H�K�F  1�H�}& Hǃ�       f���   I�FH�I�F@Hǃ�       H�KHǃ�       Hǃ       Hǃ      H�C�!  L�-�+ I�M��  H�& I�M1�fA���   I�FI��@I�^      ��       Iǅ�       Iǅ�       Iǅ       Iǅ      M�uI�E �!  H���   �   �K     H���   A��H��% H��H��- H�K8H�C    L�hH�C    L�+H�C    H�C     H�C(    H�C0    �HV��H�1+ A�����1�fD�CHH�{@H�hH�+A��H�=?% I��L�/H�O8H�G    H�G    H�G    H�G     H�G(    H�G0    ��U��A�����H�/�   fD�OHL�w@A��H�=�$ I��L�/H�O8H�G    H�G    H�G    H�G     H�G(    H�G0    �U��A�����H�/L�g@fD�WHH�='* H�O�  L�-7, E1�H��HǇ�       H�OfD���   Ƈ�    HǇ�       I�EH�I�E@HǇ�       HǇ       HǇ      H�G�s(  H�-|) H�M�  H��+ 1�Hǅ�       f���   H�Mƅ�    Hǅ�       H�PH��@Hǅ       H�U H��# Hǅ      Hǅ      H�EH�E    ��'  H�) H�K�  1�ƃ�    f���   I�EH�r# H�I�E@Hǃ�       H�KHǃ�       Hǃ�       Hǃ       Hǃ      H�C�w'  L�%�( I�L$�  H�# 1�IǄ$�       fA��$�   I�EI��@AƄ$�    I�L$IǄ$�       IǄ$�       IǄ$       IǄ$      M�l$I�$��&  �K     H���   H���   ��H�� [^_]A\A]A^�H�OH��H��, H�PH�W�  H���_��H�MH��H�{, H�PH�U�~  H����^��H�KH�_      �H�X, H�PH�S�[  H����^��I�MH��H�5, H�PI�U�8  H���^��H�OH��H�", H�PH�W�  H���^��H�MH��H��+ H�PH�U��  H���j^��H�KH��H��+ H�PH�S��  H���G^��I�L$H��H��+ H�PI�T$�  H���"^����H��(H�u% ���������tH��(�f�H�y& �����H�M& �����H�Q& �����H��& ��P��H�y& ��P��H�}& ��P���H��(�H���z�  �H��(鐚  UWVSH��(H���   L��H��H��H���Q��H��H���uR���   H������H��H��([^_]Ð������������   ����  ��Ð��������������VSH��8H�t$(H��H�A   H�A    �A  H���Q��H���   H����Q��H���Q���H��8[^Ð���UWVSH��HH�BH�AH�BH��H��H�n@H�A�B�A�B�A�B �A H�B(H�B(    H�A(H���   H��t
H9�t��  H���   H�S@H9�tFH���   H���   ���   ǃ�      ���   H���   H���   H��H[^_]�7Q���    H���   1�I�    ����ǆ�       H���   L!�H�H�
L�JH�|$8H�D$0    H�    D�D$8D�BH���   H�L$ L�L$(H��L$(�LH��H=�   u��^���WVSH��@H�AL�BL�Y@L�AL�BL�J@H�BH�AL�AD�BH�B�AD�AD�B�B�AD�AD�B �B�A D�A L�B(�B H�A(L�A(L���   H�B(H���   L9���   M9���   �@   f�L�L�L�TL�D�LD�LL�D$ L�T$(L�`      D�D$(D�DH��H=�   u�H���   H�|$8H���   H��H����N��H��H���O��H��H���O��H���uO���H��@[^_�L9�t7M9�t2L���   H���   ���   D���   D���   ���   ��     L9�t@I��I�Ѹ@   M�M� E�TE�T H��H=�   u�I���   I���   M���   �M��I��I���AUATUWVSH��   M�`E�(I�$H�\$0H��H��H�����H�@ H9���  H�CA���D$@ H�D$0H�D$8    �j  H�D$    L���  E1�1�H���I^��H�D$    L���  E1�1�H���,^��H�t$PH�VH�T$PH�H�PH9���   H�L$PH�HH�L$`H�H�@ H�L$XH��H�H�@    �� ��I��E1�1�H�D$ H����]��H�|$pH�WH�T$pH�H�PH9���   H�L$pH�HH��$�   H�H�@ H�L$xH��H�H��H�@    �yj��H�L$pH��H9�t�F�  H�L$PH��H9�t�3�  H�L$0H��H9�t� �  H��� D�mL�eH�E H�Ę   [^_]A\A]��o@)D$`�����oH)�$�   �`���H�D$    L��  E1�1�H����\������f.�     E��L��H�����w���H�L$0H��H��H9�t芐  H����W��H�L$pH��H��H9�t�l�  H��H�L$PH��H9�t�V�  H�L$0H��H9�t�C�  H���W��H����H���ȐATUWVSH��   H�t$PH��H����Y��H����I��H� H�@ H9���  H�FE1�1��D$` L�-�  H��H�D$PH�D$    H�D$X    ��[��H�H�\$0E1�L�GH�CH��H�D$0I��ba��H��������H+D$8H��a      �t  H���  A�   H���w��L�L$0H�SH�L$8L�D$XL�T$@I9�J��$  L9�H�T$PvL�VL9��  L�T$`L9���   H���2w��H�|$pH�WH�T$pH�H�PH9���   H�L$pH�HH��$�   H�H�@ H�L$xH��H�H��H�@    ��g��H�L$pH��H9�t轎  H�L$0H��H9�t誎  H�L$PH��H9�t藎  H� � �E   L�eH�E H�Đ   [^_]A\� H�L$ E1�1�H���~Z���7���f�     �o@)�$�   �K���A�   L��H�����f���A�   �����A�   �����H�t�  �>  H��H�L$0H��H9�t��  H�L$PH��H9�t���  H���HU����H����H�L$PH��H��H9�t軍  H���#U��H�L$pH��H��H9�t蝍  H��뒐�������AUATUWVSH��   M�`E�(I�$H�t$PH��H��H�t���H�@ H9���  H�FA���D$` H�D$PH�D$X    ��  H�D$    L�~�  E1�1�H���9Y��H�H�\$0E1�L�GH�CH��H�D$0I��^��H��������H+D$8H����  H�Q�  A�   H����t��L�L$0H�SH�L$8L�D$XL�T$@I9�J��G  L9�H�T$PvL�VL9��<  L�T$`L9���   H���t��H�|$pH�WH�T$pH�H�PH9���   H�L$pH�HH��$�   H�H�@ H�L$xH��H�H��H�@    �De��H�L$pH��H9�t��  H�L$0H��H9�t���  H�L$PH��H9�t��  H�T� D�mL�eH�E H�Ę   [^_]A\A]��     H�L$ E1�1�H����W���3���f�     �o@)�b      $�   �G���H�D$    L���  E1�1�H���W���S���E��L��H�����C���A�   �����A�   ����H���  ��;  H��H�L$PH��H9�t�#�  H���R��H��H�L$0H��H9�t���  ��H�L$PH��H��H9�t��  H���UR����H�L$pH��H��H9�t�͊  H��밐�������SH�� H�$� H��H��X��H��H�� [霊  ������������H��� H��X���WVSH�� H�� H��H�H�I�����H�� [^_�H��H��H����   H��H��t�Q���9�  ���������SH�� H���   H��H�� [��  ������SH��0H��� H�H��H�I�������A���~H���   �H��0[�H�T$/H������H���w   �H��0[�H��� L�A@H�H�A    L��H�A    H���   H�A    �A     H�A(    H�A0    �A8    f�H�     H���@�    H9�u�L���   H���   �A�   �D�����������������SH�� H���   H��H�� [��  ������SH�� H�� 1�H��H�����H���/���H���   H�C@H9�tH��t�ň  Hǃ�       H���   H�� [��D�����������VSH��(1�M��H�����AH��� H���A��H�CH��([^�H��H���B��H����O�����������������VSH��(1�H��H�����AH�e� H��}A��H�CH��([^�H��H���7B��H���O�����������������VSH��(1�M��H�����AH�� H��-A��H�CH��([^�H��H����A��H���?O�����������������VSH��(1�H��H�����AH�ŧ H���c      @��H�CH��([^�H��H���A��H����N�����������������SH�� H��� H�H��H�I�5A��H���]A��H��H�� [�@�  SH�� H�T� H�H��H�I�A��H��H�� [�(A����������SH�� H�$� H�H��H�I��@��H��H�� [��@����������VSH��(1�M��H�����AH�%� H���?��H�CH��([^�H��H���@��H���N�����������������VSH��(1�H��H�����AH�զ H��?��H�CH��([^�H��H���g@��H���M�����������������VSH��(1�M��H�����AH��� H��]?��H�CH��([^�H��H���@��H���oM�����������������VSH��(1�H��H�����AH�5� H��?��H�CH��([^�H��H����?��H���M�����������������SH�� H��� H�H��H�I�e?��H���?��H��H�� [�p�  SH�� H�ĥ H�H��H�I�5?��H��H�� [�X?����������SH�� H��� H�H��H�I�?��H��H�� [�(?����������SH�� H�AH��H����   H���  H�PH�CH�@    H�C�@  H�C�@H.H�C�@I,H� L� 1�A� H�S�LJH��H��$u�H�� L� 1�A� H�S�LnH��H��u�H�CH�\�  H�Z�  H�H(H�CH�@0   H�CH�P8H�CH�@@   H�� [ù�   耄  H�	� 1��@    H�H�@    H�@    �@  H�@(    H�@0    H�@8    H�@@    f�PHƀ�    H�C����������VSH��(1�M��H�QH����1҉AH�_� H������H��([^�H��H���d      �=��H���K��������������VSH��(1�M��H�A    H�����AH�� H��U����H��([^�H��H���b=��H���J������������VSH��(1�H��H�A    H����1҉AH��� H������H��([^�H��H���=��H���hJ����������VSH��(1�M��H�QH����1҉AH�o� H������H��([^�H��H����<��H���J��������������VSH��(1�M��H�A    H�����AH�� H��e����H��([^�H��H���r<��H����I������������VSH��(1�H��H�A    H����1҉AH�ˢ H������H��([^�H��H��� <��H���xI����������VSH��(H���"   H��H��([^��  H��H���ف  H���AI���VSH��(H�3 H��H��H�H�IH��tH��PH��H��([^�;��H��H���;��H����H�����������SH�� H�AH��H����   H�� H�=�  �@  H�XH�@    �@H. , L�1ҐfA�f�LPLH��H��$u�H�T L�1�fA�f��P�   H��H��u�H���  H�@0   H�X(H���  H�X8H�@@   H�� [ù�   ��  H��� �@    H�H�@    H�@    �@  H�@(    H�@0    H�@8    H�@@    �@H    ƀ�    H�C�
��������VSH��(1�M��H�QH����1҉AH�?� H�������H��([^�H��H���D:��H���G��������������VSH��(1�M��H�A    H�����AH�� H��u����H��([^�H��H����9��H���JG������������VSH��(1�H��H�A    H����1҉AH�e      �� H��#����H��([^�H��H���9��H����F����������VSH��(1�M��H�QH����1҉AH�O� H�������H��([^�H��H���T9��H���F��������������VSH��(1�M��H�A    H�����AH��� H������H��([^�H��H���9��H���ZF������������VSH��(1�H��H�A    H����1҉AH��� H��3����H��([^�H��H���8��H���F����������VSH��(H���"   H��H��([^�t~  H��H���i~  H����E���VSH��(H�� H��H��H�H�IH��tH��PH��H��([^�<8��H��H���18��H���E�����������1�H�����AH�>� H�Ð���������1�H�����AH�� H�Ð���������SH�� H�� H��H���7��H��H�� [�}  ������������H�ٞ H��7���H�ɞ H��7���1�H�����AH��� H�Ð���������1�H�����AH�ޞ H�Ð���������SH�� H�Ğ H��H��97��H��H�� [�}  ������������H��� H��7���H��� H��7���1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H��� H��H��6��H��H�� [�|  ������������H�Y� H��6���H�I� H��q6���1�H�����AH�^� H�Ð���������1�H�����AH�>� H�Ð���������SH�� H�$� H��H��6��H��H�� [��{  ������������H��� H���5���H�� H���5���SH�� H�� H��H��i  �f         H��H�� [�{  �������H�ٝ H��A  ��Q�Q �5  �����H��(	Q �QuH��(��Z�  ����������VSH��(H��H��H���|<  ��tLH���M  H���   H���a?  ��t>H����O  H���   H���>  ��t2H���O  H��   H��([^�Hǆ�       �Hǆ�       ��f�Hǆ       �А��H���   H���   ÐWVSH�� ���    H�ˉ�t���   @���   H�� [^_�D  H���   H��tQ�8 t�GYƃ�   @���   H�� [^_�@ H���x���H�H�����L�@0�    I9�tƺ    H��A�����%  ��������������VSH��(H��H���O���H���   H������1�Hǃ�       f���   1�H�����C    H���   �C H��([^Ð�����������VSH��(H��H���?���H���   H���@���H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H��([^Ð����������VSH��(H��H�������H���   H�������H���   Hǆ�       H���   ���   ���   ���   Hǃ�       ���   H��([^Ð����������VSH��(H��H������H���   H���`���H���   H���Q���H���   H���   H���   ���   H���   ���   ���   ���   ���   ���   ���   ���   H��([^Ð���������H��(H���    t�Q�Q uH��(�D  ����H�t�  �/%  ���������������ATUWVSH��0H��L��H��H���   �a3��H�t$(H��I��H������H���4��H��H���k���H���   H��tg      .L�c8H��L��� 3��H�H��H���PL��H���	4��H����3��H��H��0[^_]A\�H���H��H���3��H���3��H����>�����H��(H���   H��H���   ���҅Q�Q uH��(�H���  �<$  ������������ATUWVSH��0H9�H��H���H  ���   L�a@L�����  H�n(H��t��E1�H���y���H���   L9�tH��t�v  Hǃ�       H�������D���   H�k(E��~0E�A�1�I��I��f�H���   H�H��D�DH��I9�u��FH���   ���    D���   �CH�FH�CH�FH�CH���   H���   ��   ���    ���   ��   @���   H�|$(H���   H���r1��H���   H��H���`2��H���(2��H��H���}����   H���p����FH�ًS �C�o���H��H��0[^_]A\ÐH���   H���  �}8 ��   �}Y@���   Ɔ�   ���    �Z���H���   H����   �}8 taƃ�   �8���D  Hc�H���du  Hc��   H��H���?���H��H�     H���@�    H���u�H�n(H����������f�H������H�E H�M���H�@0H9�t��    H�����t���D  H��    �����H�E H����H�@0H9������    H���Љ������5   �����Q �8�����������H���   Ð�������VSH��(H��H������H�Ȗ H��H��H�1�Hǃ�       f���   Hǃ�       Hǃ�       Hǃ�       Hǃ       ������H��([^�H��H�������H���_;�����������������SH�� H������H�<� Hǃ�h             H�1�f���   Hǃ�       Hǃ�       Hǃ�       Hǃ       H�� [Ð��VSH��(H��H������H�ؕ H��H��H�1�Hǃ�       f���   Hǃ�       Hǃ�       Hǃ�       Hǃ       ������H��([^�H��H�������H���o:�����������������SH�� H���#���H�L� Hǃ�       H�1�f���   Hǃ�       Hǃ�       Hǃ�       Hǃ       H�� [Ð��SH�� H��� H��H��i���H��H�� [�lr  ������������H�ɔ H��A����H��� H��1�����Q�Q �  �����H��(	Q �QuH��(��
{  ����������VSH��(H��H��H���3  ��tLH��� D  H���   H���q6  ��t>H���G  H���   H���5  ��t2H���*F  H��   H��([^�Hǆ�       �Hǆ�       ��f�Hǆ       �А��H���   H���   ÐVSH��(���    H�ˉ�t���   f���   H��([^��    H���   H��t H��    �PPƃ�   f���   H��([^��  ���������������VSH��(H��H���/���H���   H�������1�ƃ�    f���   1�H�����C    Hǃ�       H���   �C H��([^Ð����VSH��(H��H������H���   H���p���H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   H��([^Ð���������VSH��(H��H������H���   H��� ���H���   Hǆ�       H���   ���   f���   ���   Hǃ�       ���   Hi      ��([^Ð���������VSH��(H��H���o���H���   H������H���   H������H���   H���   H���   ���   H���   ���   f���   ���   f���   ���   ���   ���   H��([^Ð�������H��(H���    t�Q�Q uH��(�D  ����H�T�  �  ���������������ATUWVSH��0H��L��H��H���   �A*��H�t$(H��I��H������H����*��H��H������H���   H��t.L�c8H��L��� *��H�H��H���PL��H����*��H���*��H��H��0[^_]A\�H���H��H���*��H���*��H���5�����H��(H���   H��H���   ���҅Q�Q uH��(�H�a�  �  ������������ATUWVSH��0H9�H��H���H  ���   L�a@L�����  H�n(H��t��E1�H���Y���H���   L9�tH��t�m  Hǃ�       H�������D���   H�k(E��~0E�A�1�I��I��f�H���   H�H��D�DH��I9�u��FH���   ���    D���   �CH�FH�CH�FH�CH���   H���   ��   ���    ���   ��   f���   H�|$(H���   H���R(��H���   H��H���@)��H���)��H��H�������   H���P����FH�ًS �C�o���H��H��0[^_]A\ÐH���   H����   H��    �PPƆ�   ���    ��f���   �[���H���   H��tjH��    �PPƃ�   �8���D  Hc�H���Dl  Hc��   H��H���?���H��H�     H���@�    H���u�H�n(H�����������}  �����j      ��������Q ������������H���   Ð�������VSH��(H��H�������H�(� H��H��H�1�Hǃ�       f���   ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ       �C����H��([^�H��H��� ���H���2����������SH�� H���S���H��� Hǃ�       H�1�f���   ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ       H�� [Ð�����������VSH��(H��H�������H�(� H��H��H�1�Hǃ�       f���   ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ       �C����H��([^�H��H��� ���H���1����������SH�� H���S���H��� Hǃ�       H�1�f���   ƃ�    Hǃ�       Hǃ�       Hǃ�       Hǃ       H�� [Ð�����������SH�� H�4� H��H�����H��H�� [�i  ������������H�	� H��a����H��� H��Q�����   �fi  ������Ð��������������1�H�����AH�� H�Ð���������1�H�����AH�� H�Ð���������SH�� H�ԋ H��H���"��H��H�� [��h  ������������H��� H���"���H��� H���"���1�H�����AH��� H�Ð���������1�H�����AH��� H�Ð���������SH�� H�t� H��H��i"��H��H�� [�Lh  ������������H�I� H��A"���H�9� H��1"���1�H�����AH�N� H�Ð���������1�H�����AH�.� H�Ð���������k      SH�� H�� H��H���!��H��H�� [�g  ������������H�� H��!���H�ي H��!���1�H�����AH�� H�Ð���������1�H�����AH�Ί H�Ð���������SH�� H��� H��H��I!��H��H�� [�,g  ������������H��� H��!!���H�y� H��!����   �g  ������Ð��������������H��(H�5�  H���(���������������S�|$0 A��tEI�˻�����A��D��I����D����D��E�D)�A��A��A��	G�E�w�H��L)�[�f�D�ȃ�J��@t5A�� @  I��A��҃����D��A��I�����E��A� A�u��I��D��A��I����E��A�D A�u�땐��������������S�|$0 I��tJH���������I���	fD  I��L��I��H��L��H��L��M�L)�I��	E�L E�w�H��L)�[�D�ȃ�J��@t<A�� @  I��A��H�H���I�T fD  L��I��I����M���A�u��I�ːL��I��I����M��A�D A�u�돐�S�|$0 A��tGI�˻�����A��D��I����D����D��E�D)�A��A��A��	G�HfE�w�L)�H��H��[�D�ȃ�J��@t6A�� @  I��A��҃����D��A��I�����E��A�@fA�u��I��f.�     D��A��I����E��A�D@fA�u�눐S�|$0 I��tUH���������I���	fD  I��L��I��H��L��H��L��M�L)�I��	E�L@fE�w�L)�H��H��[��    D�ȃ�J��@t:A�� @  I��A��H�H���H��L��I��I����H�M��l      A�@fA�u��I���     L��I��I����M��A�D@fA�u��|�����������������H���  H� Ð����H���  H��H�Ð�UWVS1�M�H�t$HL�T$PI�A���L��1ҐM��I)�M9�~-D�M�A��}w#M)�H9��  H��M��M�I)�M9�L���I9��  M��E1�I)�fD  B�B�	I��M9�u�J�	H��H���tQ�A�4H�h@����   D�^�1�E���L��E�
I9�D�LL�Iu�F�H��H��H��I�H�H���u�H��H���tV�A�4H�x@��~eD�^�1�E���f�     L��E�
L9�D�LL�Iu�F�H��H��H��I�H�H���u�[^_]�f.�     H��������    H���y����     H������H������ATUWVSE1�I�L�T$PH�D$X��H��1�I��I��M)�I��I9�~4D�^�A��}w*L�L)�I9��  H��I��I�M)�I��I9�H���L9��  L��H��f�H9�u�L)�H��H��H�D I�H�I��I���tWf�(A�H�p����   �K���L�\	1�fD  E�
fD�LH��L9�u��I��H��H�DI�H�I���u�H��H���tVf�(A�H�p��~f�K���L�\	1�f�     E�
fD�LH��L9�u��H��H��H�DI�H�H���u�[^_]A\�f�     I�������    H���x����     H������H�������AUATUWVSH��8H��I��1�1�M������H��H���G���H�XH���[`  I��H��H��H������H���  1��\���H�T$(H���,��H�D$(�A$H9�t�8 t:I�$    A�m      E    H��1�� ���H����_  �H��8[^_]A\A]�f.�     ���  f.�w
f.��  v�f��������  f(�fT�fU�fV��A$A�E    �H��H��t��&���db  ����AUATUWVSH��HH��I��1�1�M������H��H���7���H�XH���K_  I��H��H��H������H���  1��L���H�L$ H��L�D$8��9��H�D$8�l$ ��A�<$H9�t	�8 tA�������A�<$A�E    ���H��1������H���^  �H��H[^_]A\A]�f�     �-��  ��w�-��  ������v���������v�-��  A�<$A�E    �f.�     �-z�  ��H��H��t�%���Ea  �����AUATUWVSH��8H��I��1�1�M���b���H��H������H�XH���+^  I��H��H��H���j���H�s�  1��,���H�T$(H���?+��H�D$(�A$H9�t�8 t:A�$    A�E    H��1������H���]  �H��8[^_]A\A]�f.�     ���  .�w	.t�  v�f������a�  (�T�U�V��A$A�E    �H��H��t�$���:`  ����������H���  H� Ð����H�y�  H��H�Ð�H��t  Ð�������H��H��t  Ð����AVAUATUWVSH��0L�5P�  �   L��I��1�Ic�M�������   H��H����� ��u.L��$�   H��M��L��L�L$(�?���É�H��0[^_]A\A]A^�H���w���H�pH���\  I��H��H��H�������L��   ����M��H��L��L��$�   L�L$(�2?��H���   ���c���H���\  뉐��������AWAVAUATUWVSH��HL�l$0H��n      I��H��L��M�������|$0 ��   H�H�@�H�4H�nI9���   �~��   �� �|$$tyH��L)瀾�    ��  D���   A����D�0H�A(H�H��H�@���   H���   H�A(H;A0r�H����Ph���u�H�H�H�HًQ �������H�H�p�H�D�F E����   H�F    H�D$8H�HB��@ H��t$��  ��uH���   H��tH��P0����|  H��H��H[^_]A\A]A^A_��    H���   M��L��H��P`H�H�r�H�I9�t��V H����P���H�H�p�H�H�F    �e���f�     H�4�F ���E���H���   M��L��H��P`H�I9�H�R�H�4t�V H��������H�H�P�H�4�|$$ ������N �������L)倾�    ��   ���   @���f�@�8H�A(H�H��H�P��  H���   H�A(H;A0r�H����Ph���u�H�H�H�HًQ ���c�������H���   H��H�D$(��   H�D$(�x8 t>D�pYD���   H�Ɔ�   H�@������H�L$8H�HH�Q �������h��� L�t$(L���c���I�H�����A�    H�@0H9�t��    H�L$(��A���f�     L���   M��t`A�|$8 t)A�|$Y@���   H�Ɔ�   H�P������H�4����L������I�$H� ����    H�@0H9�t��    L���Љ���?  �:  H��H��u��Z  H�HX�K �Ct#�fa  �Z  H�H�x�H߃O �Gt"�Ha  �Ca  H���\  L���S���H������\  ����H����H���\  �א�AWAVAUATUWVSH��HL�t$0H��I��H��L�o      �M���G���|$0 ��   H�H�p�H�H�nI��I9��  �F%�   �� �D$(��   H��L)瀾�    �
  D���   A�ŉD$,�'�     fD�(H��H�A(D��f���t;H���  H���   I��H�A(H;A0r�H��T$,�PhH�H�r�H�f���I��uŋV H�������H�L�@�I�A�H ����   I�@    H�D$8H�HB��@ H��t$��  ��uH���   H��tH��P0����{  H��H��H[^_]A\A]A^A_��    H���   M��L��H��P`H�L�B�I�I9�t�A�P L�����_���H�L�@�I�I�@    �d����     �F ���I���I���   L��M��H��P`H�H�r�H�I9�I��t�V H�������H�H�p�H�I���|$( ������V �������L)倾�    ��   ���   D���#f�f�8H��H�A(��f�����   H�������H���   I��H�A(H;A0r�H�D���PhH�H�r�H�I���� H���   H����   H��    �PPf���   A��H�Ɔ�   H�p�H������D  H�L$8H�HH�Q �������i���@ H���   H��tLH��    �PPf���   ��H�Ɔ�   H�p�H�����f.�     �V H���������^����   �   H��H��u�W  H�HX�K �Ct#�]  ��V  H�H�x�H߃O �Gt"�]  �]  H����X  L�����H��������X  �f���H����H����X  �א����������H��(�   �U  H���  L�԰��H�QH��H�H�� �n]  ��������������H��8L�D$/��  H��8Ð����p      ��������H��8L�D$/��  H��8Ð������������H��(�   �2U  H���  L�$���H�QH��H�H�� ��\  ��������������H��(M�HM� �  �H��(�H��H��t�����wV  �������M� M�H��t  ����H��(�'��H��(Ð�H��(�   �T  H���  L�$���H�QH��H�H�� �^\  ��������������H��(�WX  �@����H��(Ð���������ATUWVSH��   H�t$0H�͹0   �1T  H�����H��G��I��H� H�@ H9���  H�FE1�1��D$@ L��  H��H�D$0H�D$    H�D$8    ���H�D$    L��  E1�1�H���~��H�|$PH�WH�T$PH�H�PH9��  H�L$PH�HH�L$`H�H�@ H�L$XH��H�H�@    ����I��E1�1�H�D$ H�����H�l$pH�UH�T$pH�H�PH9���   H�L$pH�HH��$�   H�H�@ H�L$xH��H�H��H�@    ��*��H�L$pH��H9�t�Q  H�L$PH��H9�t�Q  H�L$0H��H9�t�rQ  H��Y H���C   L�cH������H�K H����  L��j��H��H�x �sZ  �o@)D$`������oH)�$�   �D���A�   L��H��������H��H���V  H���\��H��H�L$0H��H9�t���P  ����H��H��H�5S H�����H�L$pH��I��H9�t�P  H�L$PH��H9�t�P  L���I���㐐������VSH��(H�ι   ��Q  H��H��H���o��L����H��H�~ �Y  H��H���NU  H�����������VSH��(H�ι   �}Q  H��H��H����q      �L�X��H��H�N �9Y  H��H����T  H���V��������H��(�'U  �@H��(Ð��������������VSH��(H�ι   �Q  H��H��H���/��L����H��H�N ��X  H��H���T  H������������VSH��(H�ι   �P  H��H��H�����L�H��H��H� �yX  H��H���>T  H�����������VSH��(H�ι   �mP  H��H��H�����L����H��H�� �)X  H��H����S  H���F��������WVSH��@H�\$ �Ϲ    �P  A��H��H��w  H���cD��H��H���'��H�L$ H��H9�t�N  H�nV H��~H�L�n��H��w  H�� H�F�W  H�L$ H��H��H9�t�AN  H���IS  H�����H���됐����������ATUWVSH�� H�YH��H�QH��M��A� H9���   �1� H)�H��~;H�I��H���P`HFH�H9���   H�H���PH���t[H�^H�VH)�H���H�W(H;W0sR�H�G(H�VH��H�^H9�sH��H�VH9�v����     H�H���PP���uPH��H�� [^_]A\�@ ��H�H���Ph���u�H��A�$ H�� [^_]A\�H�1��PH���t�H�^H�V����H�VH�^놐�������ATUWVSH�� H�AH9AH��I��L��A� ��   � 1�f���u;�   I�$L��L��H��I���P`H� H�HSH9���   H�H���PHf���t[H�SL�CI)�I���I�L$(I;L$0sLf�H��I�L$(H��H�SH;Ss^�H��H�Sf���tH�CH;Cs�� f���u�H��H�� [^_]A\���I�$L���Phf���u�Hr      ���E  H�� [^_]A\��    H�H���PP�H��PH��������������H�H� ����������H��(�   �"M  H���  L��e��H�QH��H�H� ��T  ��������������VSH��(H�ι   ��L  H��H��H���?$��L�X%��H��H�� �T  H��H���^P  H�����������VSH��(H�ι   �L  H��H��H���oo��L�p��H��H�� �IT  H��H���P  H���f��������SH�Z�I��L9�IG�1�H��tyf�     G�I���H��A8�A��H9�sE��t�A8���M���t#E��uf.�     C�I��t8�t�8����J���}wA8��!�[�f.�     E1۸   뮐�����VSH��8H�\$(H��L�D$&H������H��H��調��H�L$(�������A���~H��8[^�H�T$'H���2����H��8[^Ð���������VSH��(H�ι   �=K  H��H��H���O���L�����H��H�� ��R  H��H���N  H�����������H���  �t8������VSH��(H�ι   ��J  H��H��H������L�����H��H�� �R  H��H���^N  H�����������UVSH��H��0H�U(H��L�E0L�M8�"���H��   H  H������L�M(H)�I��H�\$ L�M�H���1 ���   �GJ  H��H��H������L����H��H���  �R  H��H����M  H��� ������������������WVSH��0H�H�P�H�\$(H��H�H��H���   ����H���@  H��H�����H�H�@�H���   H�CH9Cw�jf.�     H��H�CH9�sS� H�W0���B t0H�Cs      H�SH9�r�H�H���PP���u8H�H�H�H�Q ������H��H��0[^_��     H�H���PH���u���H�CH�S�H��H������H���#�����WVSH��0H�H�P�H�\$(H��H�H��H���   ����H���  H��H�����H�H�@�H���   H�CH9Cw'�~f.�     �H��H�Sf���tCH�CH;CsY� f���t0L�D���    H��A�Q��t.H�SH;Sr�H�H���PPf���u�H�H�H�H��Q ������H��H��0[^_�H�H���PH�H��H�����H���.����������������VSH��(H�H�@�H��H���   H��tM�{8 t�SCH������H��H��([^���� H��航��H��
   H�����H�@0H9�t�H�������������SH�� H�H�@�H��H���   H��t#H��
   �PPH��������H��H�� [� ������������������1��i������������1��i�������������;���������������K ���������������Ð��������������Ð������������SH�� H��H��y  ����H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �KO  H����H�� [Ð��������������SH�� H��H�Ay  輰��H�H��1�H9Qv)H�IH��H��tL���  E1�H�0�  ��N  H����H�� [Ð��������������SH�� H��H�y  �\���H�H��1�H9Qv)H�IH��H��tL�j�  E1�H���  �N  H����H�� [Ð��������������SH�� H��H��x  �����H�H��1�H9Qv)H�IH��H��tL�*�  E1�H�p�  �+N  H��t      ��H�� [Ð��������������SH�� H��H�ax  蜯��H�H��1�H9Qv)H�IH��H��tL���  E1�H��  ��M  H����H�� [Ð��������������SH�� H��H�x  �<���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �kM  H����H�� [Ð��������������SH�� H��H��w  �ܮ��H�H��1�H9Qv)H�IH��H��tL���  E1�H�P�  �M  H����H�� [Ð��������������SH�� H��H�qw  �|���H�H��1�H9Qv)H�IH��H��tL�j�  E1�H���  �L  H����H�� [Ð��������������SH�� H��H�!w  ����H�H��1�H9Qv)H�IH��H��tL�*�  E1�H���  �KL  H����H�� [Ð��������������SH�� H��H��v  輭��H�H��1�H9Qv)H�IH��H��tL�
�  E1�H�0�  ��K  H����H�� [Ð��������������SH�� H��H��v  �\���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �K  H����H�� [Ð��������������SH�� H��H�1v  �����H�H��1�H9Qv)H�IH��H��tL���  E1�H�p�  �+K  H����H�� [Ð��������������SH�� H��H��u  蜬��H�H��1�H9Qv)H�IH��H��tL�j�  E1�H��  ��J  H����H�� [Ð��������������SH�� H��H��u  �<���H�H��1�H9Qv)H�IH��H��tL�*�  E1�H���  �kJ  H����H�� [Ð��������������SH�� H��H��p  �ܫ��H�H��1�H9Qu      v)H�IH��H��tL�
�  E1�H�P�  �J  H����H�� [Ð��������������SH�� H��H�qp  �|���H�H��1�H9Qv)H�IH��H��tL�*�  E1�H���  �I  H����H�� [Ð��������������SH�� H��H�1p  ����H�H��1�H9Qv)H�IH��H��tL�J�  E1�H���  �KI  H����H�� [Ð��������������SH�� H��H��o  輪��H�H��1�H9Qv)H�IH��H��tL�
�  E1�H�0�  ��H  H����H�� [Ð��������������SH�� H��H�q�  �\���H�H��1�H9Qv)H�IH��H��tL�Z�  E1�H���  �H  H����H�� [Ð��������������SH�� H��H�!�  �����H�H��1�H9Qv)H�IH��H��tL�:�  E1�H�p�  �+H  H����H�� [Ð��������������SH�� H��H�A�  蜩��H�H��1�H9Qv)H�IH��H��tL�:�  E1�H��  ��G  H����H�� [Ð��������������SH�� H��H���  �<���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �kG  H����H�� [Ð��������������SH�� H��H��r  �ܨ��H�H��1�H9Qv)H�IH��H��tL���  E1�H�P�  �G  H����H�� [Ð��������������SH�� H��H�1r  �|���H�H��1�H9Qv)H�IH��H��tL�z�  E1�H���  �F  H����H�� [Ð��������������SH�� H��H��q  ����H�H��1�H9Qv)H�IH��H��tL�:�  E1�H���  �KF  H����H�� [Ð������v      ��������SH�� H��H��q  輧��H�H��1�H9Qv)H�IH��H��tL���  E1�H�0�  ��E  H����H�� [Ð��������������SH�� H��H�Aq  �\���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �E  H����H�� [Ð��������������SH�� H��H��p  �����H�H��1�H9Qv)H�IH��H��tL�z�  E1�H�p�  �+E  H����H�� [Ð��������������SH�� H��H��p  蜦��H�H��1�H9Qv)H�IH��H��tL�j�  E1�H��  ��D  H����H�� [Ð��������������SH�� H��H�qp  �<���H�H��1�H9Qv)H�IH��H��tL�J�  E1�H���  �kD  H����H�� [Ð��������������SH�� H��H�!p  �ܥ��H�H��1�H9Qv)H�IH��H��tL�*�  E1�H�P�  �D  H����H�� [Ð��������������SH�� H��H��o  �|���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �C  H����H�� [Ð��������������SH�� H��H��o  ����H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �KC  H����H�� [Ð��������������SH�� H��H�1o  輤��H�H��1�H9Qv)H�IH��H��tL���  E1�H�0�  ��B  H����H�� [Ð��������������SH�� H��H��n  �\���H�H��1�H9Qv)H�IH��H��tL�j�  E1�H���  �B  H����H�� [Ð��������������SH�� H��H��n  �����H�H��1�H9Qv)H�IH��H��tLw      �*�  E1�H�p�  �+B  H����H�� [Ð��������������SH�� H��H�An  蜣��H�H��1�H9Qv)H�IH��H��tL�Z�  E1�H��  ��A  H����H�� [Ð��������������SH�� H��H��m  �<���H�H��1�H9Qv)H�IH��H��tL��  E1�H���  �kA  H����H�� [Ð��������������SH�� H��H��m  �ܢ��H�H��1�H9Qv)H�IH��H��tL���  E1�H�P�  �A  H����H�� [Ð��������������SH�� H��H�Qm  �|���H�H��1�H9Qv)H�IH��H��tL���  E1�H���  �@  H����H�� [Ð��������������H��(H���  H��m����������������SH�� H��H�aj  �����H�H9BH�Jv*H��H��t!L���  E1�H�u�  �0@  H��tH�� [��������7  �����������SH�� H��H�j  蜡��H�H9BH�Jv*H��H��t!L�o�  E1�H��  ��?  H��tH�� [��`����{7  �����������SH�� H��H��i  �<���H�H9BH�Jv*H��H��t!L�O�  E1�H���  �p?  H��tH�� [�� ����7  �����������SH�� H��H�qi  �ܠ��H�H9BH�Jv*H��H��t!L�/�  E1�H�U�  �?  H��tH�� [������6  �����������SH�� H��H�!i  �|���H�H9BH�Jv*H��H��t!L���  E1�H���  �>  H��tH�� [��@����[6  �����������SH�� H��H��h  ����H�H9BH�Jv*H��H��t!L�O�  E1�H���  �P>  H��tH��x       [��������5  �����������SH�� H��H��h  輟��H�H9BH�Jv*H��H��t!L��  E1�H�5�  ��=  H��tH�� [������5  �����������SH�� H��H�1h  �\���H�H9BH�Jv*H��H��t!L���  E1�H���  �=  H��tH�� [�� ����;5  �����������SH�� H��H��g  �����H�H9BH�Jv*H��H��t!L���  E1�H�u�  �0=  H��tH�� [��������4  �����������SH�� H��H��g  蜞��H�H9BH�Jv*H��H��t!L���  E1�H��  ��<  H��tH�� [��`����{4  �����������SH�� H��H�Ag  �<���H�H9BH�Jv*H��H��t!L�O�  E1�H���  �p<  H��tH�� [�� ����4  �����������SH�� H��H��f  �ܝ��H�H9BH�Jv*H��H��t!L�/�  E1�H�U�  �<  H��tH�� [������3  �����������SH�� H��H��f  �|���H�H9BH�Jv*H��H��t!L��  E1�H���  �;  H��tH�� [��@����[3  �����������SH�� H��H�Qf  ����H�H9BH�Jv*H��H��t!L���  E1�H���  �P;  H��tH�� [��������2  �����������SH�� H��H�f  輜��H�H9BH�Jv*H��H��t!L���  E1�H�5�  ��:  H��tH�� [������2  �����������SH�� H��H��e  �\���H�H9BH�Jv*H��H��t!L�O�  E1�H���  �:  H��tH�� [�� ����;2  �����������SH�� H��H��`  �����H�H9BH�Jvy      *H��H��t!L�/�  E1�H�u�  �0:  H��tH�� [��������1  �����������SH�� H��H��`  蜛��H�H9BH�Jv*H��H��t!L��  E1�H��  ��9  H��tH�� [��`����{1  �����������SH�� H��H�1`  �<���H�H9BH�Jv*H��H��t!L���  E1�H���  �p9  H��tH�� [�� ����1  �����������SH�� H��H��_  �ܚ��H�H9BH�Jv*H��H��t!L���  E1�H�U�  �9  H��tH�� [������0  �����������SH�� H��H��_  �|���H�H9BH�Jv*H��H��t!L���  E1�H���  �8  H��tH�� [��@����[0  �����������SH�� H��H�A_  ����H�H9BH�Jv*H��H��t!L�o�  E1�H���  �P8  H��tH�� [��������/  �����������SH�� H��H�Ѻ  輙��H�H9BH�Jv*H��H��t!L���  E1�H�5�  ��7  H��tH�� [������/  �����������SH�� H��H���  �\���H�H9BH�Jv*H��H��t!L���  E1�H���  �7  H��tH�� [�� ����;/  �����������SH�� H��H���  �����H�H9BH�Jv*H��H��t!L���  E1�H�u�  �07  H��tH�� [��������.  �����������SH�� H��H�Q�  蜘��H�H9BH�Jv*H��H��t!L�_�  E1�H��  ��6  H��tH�� [��`����{.  �����������SH�� H��H��a  �<���H�H9BH�Jv*H��H��t!L��  E1�H���  �p6  H��tH�� [�� ����.  ���z      ��������SH�� H��H��a  �ܗ��H�H9BH�Jv*H��H��t!L���  E1�H�U�  �6  H��tH�� [������-  �����������SH�� H��H�Aa  �|���H�H9BH�Jv*H��H��t!L���  E1�H���  �5  H��tH�� [��@����[-  �����������SH�� H��H��`  ����H�H9BH�Jv*H��H��t!L�_�  E1�H���  �P5  H��tH�� [��������,  �����������SH�� H��H��`  輖��H�H9BH�Jv*H��H��t!L��  E1�H�5�  ��4  H��tH�� [������,  �����������SH�� H��H�Q`  �\���H�H9BH�Jv*H��H��t!L���  E1�H���  �4  H��tH�� [�� ����;,  �����������SH�� H��H�!`  �����H�H9BH�Jv*H��H��t!L���  E1�H�u�  �04  H��tH�� [��������+  �����������SH�� H��H��_  蜕��H�H9BH�Jv*H��H��t!L���  E1�H��  ��3  H��tH�� [��`����{+  �����������SH�� H��H��_  �<���H�H9BH�Jv*H��H��t!L���  E1�H���  �p3  H��tH�� [�� ����+  �����������SH�� H��H�1_  �ܔ��H�H9BH�Jv*H��H��t!L�O�  E1�H�U�  �3  H��tH�� [������*  �����������SH�� H��H��^  �|���H�H9BH�Jv*H��H��t!L��  E1�H���  �2  H��tH�� [��@����[*  �����������SH�� H��H��^  ����H�H9BH�Jv*H��H��t!L��� {       E1�H���  �P2  H��tH�� [��������)  �����������SH�� H��H�A^  輓��H�H9BH�Jv*H��H��t!L���  E1�H�5�  ��1  H��tH�� [������)  �����������SH�� H��H��]  �\���H�H9BH�Jv*H��H��t!L���  E1�H���  �1  H��tH�� [�� ����;)  �����������SH�� H��H��]  �����H�H9BH�Jv*H��H��t!L���  E1�H�u�  �01  H��tH�� [��������(  �����������SH�� H��H�Q]  蜒��H�H9BH�Jv*H��H��t!L��  E1�H��  ��0  H��tH�� [��`����{(  �����������SH�� H��H�]  �<���H�H9BH�Jv*H��H��t!L�?�  E1�H���  �p0  H��tH�� [�� ����(  �����������SH�� H��H��\  �ܑ��H�H9BH�Jv*H��H��t!L���  E1�H�U�  �0  H��tH�� [������'  �����������VSH��(H��H��H��t H���ה��H��H��I������H��H��([^�H�H�H�H�Q ���Z���H��H��([^�VSH��(H��H��H��t H��臔��H��H��I���i���H��H��([^�H�H�H�H�Q ���
���H��H��([^�VSH��(H��H��H��t H���7���H��H��I������H��H��([^�H�H�H�H�Q ��躬��H��H��([^�H��8A�   �T$/H�T$/�����H��8Ð��H��(A�   �T$8H�T$8����H��(Ð��H��8A�   �T$/H�T$/����H��8Ð��H��H�	L�A�I�A	PÐ�������������H��H�	Hc�H�I�H�TÐ����|      ��������H��H�	��L�A�I�A!PÐ�����������H��H�	Hc�H�I�H�TÐ������������H��H�	L�A�@   I���t��
�   t1Ƀ�����A�P��	�A�PÐ�����UWVSH��(H�H�p�H�ˉ�H΀��    tH��@���   H��([^_]�H���   H��t9�}8 tƆ�   ��f�H��訇��H�E H�݉��H�@0H9�tٺ    H�������������VSH��(H��H��H��t H������H��H��I������H��H��([^�H�H�H�H�Q ������H��H��([^�AUATUWVSH��(H��H��H����   H������I��H��������?I9���   K�,$H����"  M��I��taH��H�@�H���   H����   I�l-�L��H���*f.�     H�H��H���V�H�@�H���   H��tYH��PPH9�f�u�M��L��H���4���L���<"  H��H��([^_]A\A]�H�H�H�H��Q �������H��H��([^_]A\A]�����H��H��u6�D$  H�Hx�O �Gt>��*  �+  H��H��L����!  H��H�����$  H�H�p�H��N �Ft�*  �*  H���&  H��������%  �J���H����%  H�������������H��(A�   f�T$8H�T$8�G���H��(Ð�H��H�	L�A�I�A	PÐ�������������H��H�	Hc�H�I�H�TÐ������������H��H�	��L�A�I�A!PÐ�����������H��H�	Hc�H�I�H�TÐ������������H��H�	L�A�@   I���t��
�   t1Ƀ�����A�P��	�A�PÐ�����WVSH�� H�H�p�H�ˉ�H΀��    tH��f���   H�� [^_}      �H���   H��tH��    �PPƆ�   �����������������SH��0H�H�@�H����H���   H��t$H��PPH�T$.A�   H��f�D$.�����H��0[�������������ATUWVSH�� H��L��H��L�cH���ю��L�#H��H�C    H���C H�WH��0��H��������H+CH9�w+I��H��H�����L�GH��H����H��H�� [^_]A\�H�q  �����H�H��I9�t�V  H��������������������WVSH�� E1�H�yL��H��H�9H�L�BH��I������L�FH��H����H��H�� [^_�H�H��H9�t��  H���U��������UWVSH��8H�i�A ��H��H�)L��H�A    I�@H�P�0��H�S@��E1�H�ى|$ A�   ����L�FH��H����H��H��8[^_]�H�H��H9�t�h  H�����������������������ATUWVSH��0H��H��L��L�d$/H���0���1�1�M��H���A���H��H�H�H�P�H�����I��H��H���ޙ��H��H���Ú��H��H��0[^_]A\�H�H��L��H������H���;��������������VSH��8H�L��D�@�H��H�H�H�QE��x ��H�H��H���^���H��H��8[^�@ H�T$/E1��c�����H�H�T$/H��H��蝕��H������������UWVSH��8H�|$/H��L��1ɉ�I��1��O���H��H�H�H�P�H������D�ź   H���H���H��H���͙��H��H��8[^_]�H�H��H��H������H���G����������ATUWVSH�� H��L��H��L�cH���Y���H�C    H�WH��H��1�L�#f�CH��n,��H��������?H+CH9�w+I��~      H��H����-��L�GH��H���-��H��H�� [^_]A\�H�wq  �����H�H��I9�t�4  H������������������WVSH�� E1�H�yL��H��H�9H�H�RL�PH������L�FH��H��g-��H��H�� [^_�H�H��H9�t��  H���4�������UWVSH��81�H�A    ��H��L��f�AI�@H�iH�)H�P�n+��H�S��A�   E1��|$ H���R��L�FH��H���,��H��H��8[^_]�H�H��H9�t�G  H���������������������ATUWVSH��0H��H��L��L�d$/H��踉��1�1�M��H���q��1�H��f�PH���@�    H�@�    H�H�H�P�H��� ��I��H��H������H��H�����H��H��0[^_]A\�H�H��L��H������H��������VSH��8H�L��D�@�H��H�H�H�QE��x ��H�H��H���^��H��H��8[^�@ H�T$/E1��3����H�H�T$/H��H���]��H�����������UWVSH��8H�|$/H��L��1ɉ�I��1��o��1�H��f�PH���@�    H�@�    H�H�H�P�H������D�ź   H���?��H��H�����H��H��8[^_]�H�H��H��H������H����������������������;   ������������+   ������������K  ������������;  �����������AWAVAUATUWVSH��HE1�H��H��H�L$7H����V���|$7 H�E �?  H�P�H�\$8H��������H��H�L�bM��LN�H���   �K���H������H��I������H�E H�@�H���   H�CH9C��  � M�l$�1�L9���   �����  M�N0��A�Q �      �   L�CL��H�SH)�H��M��I)�L9�IO�H����   H�BH�H9���   D�RC�Q t��   f�D�C�Q u	H��H9�w�I��I)�M����   L�L�L9�H�C��   L9�� �W�������  � H�E H��H�P�H�D    u�   H�H�H�Q �h���H��H��H[^_]A\A]A^A_�@ �H�CL�H��H�SH9�siH��H�CH9���   � L�������A�   A�   M��H��L�L$(L�辆��L�L$(H�CL�CL�L�L9�H�C�4���H�H���PH����H�H���PP���uJA� H�E H��H�P�H�D    ҃����%���H�H���PH�7���H�H���PHL���-���I���H�CH�S�:���H��H��u8��  H�E Hh�M �Etl�  1���H��H��H�������H��H��1���  H�E H�x�H�O �Gt�K  �  H�������H�E �   �x���H���  H�������  H���  H����������������VSH��8E1�H��H��H�L$/H���S���|$/ t&H�H�@�H���   H�AH9Av�H��H�A�H��H��8[^�H��PP���uH�H�H�HًQ ���M���H��H��8[^É��H��H��u�  H�HX�K �Ct#�Y  �  H�H�p�HރN �Ft�;  �6  H���  H�������  �e���H���  H������������������H��H�	L�A�I�A	PÐ�������������H��H�	Hc�H�I�H�TÐ������������H��H�	��L�A�I�A!PÐ�����������H��H�	Hc�H�I�H�TÐ������������H��H�	L��      A�@   I���t��
�   t1Ƀ�����A�P��	�A�PÐ�����UWVSH��(H�H�p�H�ˉ�H΀��    tH��@���   H��([^_]�H���   H��t9�}8 tƆ�   ��f�H���x��H�E H�Mz��H�@0H9�tٺ    H�������s������AVAUATUWVSH��0E1�I��H��H�L$'L�������|$' I�$��   H�P�H�\$(H��������H��L�H�zH��HN�H���   �����H������H��H������I�$H�@�I���   H�CH9C�  D�0L�l~�1�L9�tefA����  H�E E�ƺ    H���P����   H��H��H�SfD�v�H;Ss�H��H�Sf���t}H�CH;C��   L9�D�0u�fA�����   I�$1�H��fA�U H�P�I�D    u�   H�H�L�Q �[���L��H��0[^_]A\A]A^�f�     H�H���PPf���u�I�$f�  H�P�I�D    �   �@ H�H���PHA�������H�H���PHA�������I���Z���1�H��f�I�$H�P�I�D    ҃����U���H��H��u<�!  I�$L`�A�L$ A�D$tl�  1���H��H��H�������H��H��1����  I�$H�H�L�I �At�{  ��  H�������I�$�   �����H����  H��������J  H���  H����������������VSH��8E1�H��H��H�L$/H��蔵���|$/ t-H�H�@�H���   H�QH9Qv$�H��H�Qf���t#f�H��H��8[^�fD  H��PP���     H�H�H�HًQ ��苡��H��H��8[^�H��H��u��  H�HX�K �Ct#�}�        ��  H�H�p�HރN �Ft�_  �Z  H����  H��������  �`���H���  H����������������������H��H�	L�A�I�A	PÐ�������������H��H�	Hc�H�I�H�TÐ������������H��H�	��L�A�I�A!PÐ�����������H��H�	Hc�H�I�H�TÐ������������H��H�	L�A�@   I���t��
�   t1Ƀ�����A�P��	�A�PÐ�����WVSH�� H�H�p�H�ˉ�H΀��    tH��f���   H�� [^_�H���   H��tH��    �PPƆ�   ��躺������������SH�� H��  H�H���  H��H�A�H�̣  H�IH�A�    H��H��ą��H�K�H�� [��  ������H���  H�H�G�  H��H�A�H���  H�A�    H��H��|���������������VSH��(H�� H�A�H�q�H��PH��H���   H�IH��(H�A�H�� H��20��H�KP�y���H��  H�K@H��H�C�a���H�"�  H�C�    H�H���  H�C�H�ݢ  H���   H��H���   �ք��H��H��([^��  ��������SH�� H�L H�A�H��PH��H���   H�IH��(H�A�H� H��/��H�KP�����H�7�  H�K@H��H�C����H�w�  H�C�    H�H��  H�C�H�2�  H���   H��H���   H�� [�&���������VSH��(H�+ H�A�H�q�H��PH��H���   H�IH��(H�A�H�� H��BR��H�KP�)���H���  H�K@H��H�C����H��  H�C�    H�H��  H�C�H���  H���   H��H���   膃�      ��H��H��([^�  ��������SH�� H�| H�A�H��PH��H���   H�IH��(H�A�H�O H��Q��H�KP�~���H���  H�K@H��H�C�f���H�G�  H�C�    H�H�e�  H�C�H��  H���   H��H���   H�� [�ւ��������SH�� H�<�  H�H��  H��H�A�H���  H�IH�A�    H��H�蔂��H�K�H�� [�  ������H��  H�H���  H��H�A�H�`�  H�A�    H��H��L���������������SH�� H�H�X�H�%�  H�H�CH�Ǫ  H�H��  H�KH�C    H��H�C�����H��H�� [��
  ���������������H�HH�H�ʪ  H�AH�o�  H��H�A�H���  H�A�    H��H�餁������SH�� H�H�X�H�� H�H�H�p�  H�KH�C    H��H�C�g���H��H�� [�j
  ����������H�HH�H�� H�H�(�  H��H�A�    H��H�� ���SH�� H�H�X�H�� H�H�H��  H�KH��H�C����H��H�� [��	  ��H�HH�H�� H�H���  H��H��H�鸀����������SH�� H�H�X�H�5 H�H�H�KH��PH���   H��(H�CH�	 H�C�p+��H�K`����H� �  H�KPH��H�C����H�`�  H�C    H�CH���  H�H��  H���   H��H���   ����H��H�� [�	  �������SH�� H�H�X�H�� H�H�H�KH��PH���   H��(H�CH�Y H�C��*��H�K`����H�p�  H�KPH��H�C�����H���  H�C    �      H�CH�M�  H�H�k�  H���   H��H���   H�� [�_�����������������SH�� H�H�X�H�U H�H�H�KH��PH���   H��(H�CH�) H�C�pM��H�K`�W���H�К  H�KPH��H�C�?���H� �  H�C    H�CH�=�  H�H�˜  H���   H��H���   �~��H��H�� [�  �������SH�� H�H�X�H�� H�H�H�KH��PH���   H��(H�CH�y H�C��L��H�K`����H� �  H�KPH��H�C����H�p�  H�C    H�CH���  H�H��  H���   H��H���   H�� [��}�����������������SH�� H�H�X�H�u H�H�H�Л  H�KH�C    H��H�C�}��H��H�� [�  ����������H�HH�H�* H�H���  H��H�A�    H��H��p}��SH�� H�H�X�H�E H�H�H�P�  H�KH��H�C�?}��H��H�� [�B  ��H�HH�H�
 H�H��  H��H��H��}����������SH�� H�H�X�H�U H�H�H�KH��(H���   H�a H�C��'��H�KX����H�x�  H�KHH��H�C�����H�(�  H�C    H�H�~�  H���   H��H���   �w|��H��H�� [�z  ����������SH�� H�H�X�H�� H�H�H�KH��(H���   H�� H�C�('��H�KX�o���H�ؗ  H�KHH��H�C�W���H���  H�C    H�H�ޙ  H���   H��H���   H�� [��{����SH�� H�H�X�H�u H�H�H�KH��(H���   H�� H�C��I���      H�KX�����H�X�  H�KHH��H�C�����H�H�  H�C    H�H�^�  H���   H��H���   �G{��H��H�� [�J  ����������SH�� H�H�X�H�� H�H�H�KH��(H���   H� H�C�XI��H�KX�?���H���  H�KHH��H�C�'���H���  H�C    H�H���  H���   H��H���   H�� [�z����SH�� H�H�X�H��  H�H�CH���  H�H�u�  H�KH�C    H��H�C�\z��H��H�� [�_  ���������������H�HH�H���  H�AH�O�  H��H�A�H��  H�A�    H��H��z������SH�� H�H�X�H�u H�H�H�KH��(H���   H�a H�C��$��H�KP����H�x�  H�K@H��H�C�����H�h�  H�H���  H���   H��H���   �y��H��H�� [�  ��SH�� H�H�X�H�� H�H�H�KH��(H���   H��
 H�C�8$��H�KP����H��  H�K@H��H�C�g���H�إ  H�H���  H���   H��H���   H�� [��x������������SH�� H�H�X�H�� H�H�H�KH��(H���   H��
 H�C�G��H�KP�����H�h�  H�K@H��H�C�׽��H���  H�H�v�  H���   H��H���   �_x��H��H�� [�b  ��SH�� H�H�X�H� H�H�H�KH��(H���   H�1
 H�C�xF��H�KP�_���H�ؓ  H�K@H��H�C�G���H��  H�H��  H���   H��H���   H�� [��w������������SH�� H��H�	�AX    Ɓ�    ���H��      1�f�PyH�PhH�@(    H�@     H�@0    H�PH�PH�P�P\�P`�PdH�� [Ð�SH�� H��H�	�AX    Ɓ�    �A��H�1�f�PyH�PhH�@(    H�@     H�@0    H�PH�PH�P�P\�P`�PdH�� [Ð��   �������������o������������������������������   ������������{   �����������SH�� �   H��H��HD�H���,o��H��tH�� [�f�     �{���H��t���ֹ   ��   H�A�  L�ʃ��H��H��H�H�i�  �  ����VSH��(�   H��H��HD�H���n��H��H��tH��H��([^Ð����H��t�����H��t�w���H���?  �Z  �͐�������WH�� ��   �in��H��H��t1�H�׹   �H�H��H�� _� ��   �f���H��H��u��������������WSH��(H���   H���n��H��H��t#1�H�׹   �H�H���   H��([_��     H������H��H��u����������������H��(�   ����H���  L��Z��H�QH��H�H�s�  �N  ��������������H��(�   �R���H�k�  L�Ԓ��H�QH��H�H���  �  ��������������SH�� H���  L�C�H� �Լ����HH�H��vH��uKL� 1�H�� [�f�     D�Sغ   D)�E��A��A�RAHщS؃hL9�tH�K�L� H�C�H�� [���������SH�� H��H��t�n���H� �Լ����HH��v����H�K�������������������ATUWVSH��PH���.���H�C�H�K�H�k�Hcs�H�{�H�D$0� ���H�������#  H� �@PL����         uMH�\$ H��1�I������I��$p���I��M��H��������u;I��E1�H��H�ײ  �һ����u'H���V���L� �H���   �   H�������7  �   ����H�V�  L���H��H��H�H�~�  �Y  ���������H��(�W  H�H��t�BPH�tH��p���H��(�f.�     1�H��(Ð��������H��(A�   �   H�ZS  ��k��� �������������������H��(��   H�H��t%H� �Լ����HQPH��w+�Q(��x��t3xE�Q(H��(�D  ��u�L�A L� ��f�H��PH�     H��(����H�Q H��PH�H��(�����������H��  H9�vH�  H9�s�S��� ��j�������������H��  H��   H9�vH�  H9�s�����j���������H�A�Ð����������H��:  ������������������������VSH��(H�S���H��H�:  �4���H�m#  ��}����um�C H�	���H��9  ����H�6#  �Av����uAH�6#  �1�����uH��([^�H�5�  �   �u���L�����H�0H��  H���<  �w����B���H��H����  H��H��H��u
�����H�����<���������������AUATUWVSH��(E1����H��tD��H��([^_]A\A]��    H�Y���H�"9  �=���H�v"  ��|����A����   H�=���H�-�8  L�%!����:�{ tyH��H�������L��H�5$"  H��8  ����H�!"  H���9v����ue�; t�H�	"  ������U���H�=��  �   �K���L�����H�8H���  H���  f�H��!  �CA�  �       �~���������H�=y�  �   �����L�(���H�8H�N�  H����  �����H���Y  H�������VSH��(H�3���H��H��7  ����H�M!  �{����up�C H�����H��7  �����H�!  �t����uAH�!  �~����uH��([^�H�5��  �   �R���L�����H�0H���  H���  �T�������H��H���  H��H��H��u
����H�����������������SH�� ǁ`���    H��H��p���L��x����K���H�C��ғ��H�C�H� ++CCUNGH�C�H�����H�C�H��`���H�� [Ð�������H��(A�   �   H��N  �]g����������������������SH�� �V���H��@H��t/H� �Լ����HQPH��v H�     H�YPH������H�������6����Y(��WVSH�� H��H��L�������H��@�@�C�    H�{�H�s��_���H�C������C�   H�C�H� ++CCUNGH�H�����H�CH���{���H������辿����������������H��(�   ����H���  L�t���H�QH��H�H�Ӳ  �N�����������������UWVSH��hH�H��H�P�H��L��L��H�H�H�H�       H�D$@    H�D$PH�H�D$H    H9H�utH�L�D$@H�T$ I��L�D$8H��A�   H�\$0H�l$(�P8L�D$@M��L��t<D�L$PD�ʃ���t.�T$L�L$H!у���t����tE��uH��xL�H9�t71�H��h[^_]�D  H���t�H�H�\$ I��H��H���P@����u�L�D$@L��H��h[^_]Ð������������H��8H�%���H�D$ ����H��8Ð�����H��4  �      T|������H�I4  �D|������H�I  �4|������H�I�  H�B4  H�;4  鶀��������Ð��������������Ð���������������=�   u��  �=�   u��  �=�   u��  �=�   u��  �=)   u�   �=9   u�0  �=�   u��  �=�   u��  Ð���������������=y   u�p  �=y   u�p  �=	   u�   �=   u�  �=�   u��  �=�   u��  �=i   u�`  �=9   u�0  Ð���������������=i   u�`  �=i   u�`  �=�   u��  �=�   u��  �=	   u�   �=�   u��  �=�   u��  �=9   u�0  �=	   u�   �=�   u��  �=�   u��  �=   u�  Ð���������������=�   u��  �=�   u��  �=�   u��  �=�   u��  �=I   u�@  �=�   u��  �=�   u��  �=y   u�p  �=I   u�@  �=   u�  �=�   u��  �=Y   u�P  Ð��������������H��(H�5
  1���x��� $ H�6
   $ �a��H��H�
  t&H�
  H�  $ H�@    H�����H��(���H��	      H��	      �ؐ��������������H��(H�  �w����t+�   �b���H���  H�L�����H��H�ǖ  �"����H��(Ð������������      H��(H�E����0��H�I���H��(� ��H�D$(    H�%   H�D$(    H�%   �%        H�D$(    H�%   H�D$(    H�%   H�D$(    H�%   H�D$(    H�%   H�D$(    H�%   H�D$(    H�%   �����������VSH��8H�D$XH�˹   H�T$XL�D$`L�L$hH�D$(�`��A�   �   H��m  I���z_��H�t$(�   �`��H��H��I���]^����_���������������������������������@     g@     @
J     �
J     `J     0J      J     �J     J             ��������                                                                                                                                
               �J             ��������        ����            �                              5   �����                       k���h                     ����            @   ÿ���?                    ��L             �oA             �oA     �oA     �oA             �oA             ��������        ����������������������������    �����������������J             �J             �J             �J             �J             �J             ��J     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��A             �I                                                                                                                                                                                                                                                                                                             �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��J             ��J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                      �XJ             �XJ             YJ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �YJ     �      �YJ                     YJ     $YJ     ,YJ     6YJ     >YJ     FYJ     NYJ     VYJ     ^YJ     fYJ     nYJ     vYJ     FYJ     ~YJ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                      P�J                                                                                                           2��-�+          �] �f���                                                                                                                                                                                                                                                                                                         hello world!                   __gnu_cxx::__concurrence_lock_error     __gnu_cxx::__concurrence_unlock_error basic_string::append      locale::_S_normalize_category category not found        locale::_Impl::_M_replace_facet __gnu_cxx::__concurrence_lock_error     __gnu_cxx::__concurrence_unlock_error *                                  true false t r u e   f �      a l s e                  true false t r u e   f a l s e                 uninitialized __any_string  ����t���t���t���t���t���t���t���t������t���t���t���t���t���t���4���t���t���4���t���t���|���<���<���<���<���<���<���<���<�������<���<���<���<���<���<�������<���<�������<���<���    cannot create shim for unknown locale::facet    %s: __pos (which is %zu) > this->size() (which is %zu)  basic_string::at: __n (which is %zu) >= this->size() (which is %zu) basic_string::copy basic_string::compare basic_string::_S_create basic_string::erase basic_string::_M_replace_aux basic_string::insert basic_string::replace basic_string::assign basic_string::append basic_string::resize basic_string::_S_construct null not valid basic_string::basic_string basic_string::substr /dev/urandom default /dev/random      random_device::random_device(const std::string&) rb mt19937             %s: __pos (which is %zu) > this->size() (which is %zu)  basic_string::at: __n (which is %zu) >= this->size() (which is %zu) basic_string::copy b�      asic_string::compare basic_string::_S_create basic_string::erase basic_string::_M_replace_aux basic_string::insert basic_string::replace basic_string::assign basic_string::append basic_string::resize basic_string::_S_construct null not valid basic_string::basic_string basic_string::substr               C POSIX         C POSIX space print cntrl upper lower alpha digit punct xdigit alnum graph blank                basic_string::append C POSIX basic_string::erase        %s: __pos (which is %zu) > this->size() (which is %zu)  �D��`D��1D��D���D��l<���;���;���;���<��%.*Lf %m/%d/%y %H:%M %H:%M:%S   ����x������������������:���8���������������������������؏������h�����������������������������������������8���8���(���h���8���������8���������������(����������������������x�������������������D���t��D����D���@���p���@��� ���@���            uninitialized __any_string  $���������������������������d�������������������������������������������������������������      ����������������,���������������������������l�����������l�����������    cannot create shim for unknown locale::facet    basic_string::append C POSIX basic_string::erase        %s: __pos (which is %zu) > this->size() (which is %zu)  �U��0U���T��sT���U���L��\L��L���K���L��%.*Lf %m/%d/%y %H:%M %H:%M:%S   ��������x���X�������������������x��������������������������������������������������������������x���Y�����������������������������������x�������������������������������������������z�����������������������X������������������x��� ��2#���!���!��J ��\��n����������            basic_filebuf::underflow codecvt::max_length() is not valid     basic_filebuf::underflow invalid byte sequence in file  basic_filebuf::underflow incomplete character in file   basic_filebuf::underflow error reading the file basic_filebuf::xsgetn error reading the file    basic_filebuf::_M_convert_to_external conversion error          basic_ios::clear                ios_base::_M_grow_words allocation failed       ios_base::_M_gro�      w_words is not valid            C POSIX basic_string::erase     %s: __pos (which is %zu) > this->size() (which is %zu)  x���X���8������������������d���D�������%.*Lf %m/%d/%y %H:%M %H:%M:%S   ��������������� ��� ��� ���B���p��� ��� ��� ���C��� ��� ��� ��� ������p���@��� ��� ��� �������������� ��� ��� ��� ��� ��� ���@���@���0���c���0��� ��� ���@��� ��� ��� ��� ��� ������� ��� ��� ��� ��� ���P��� ��� ��� �����������S��lV��|U��lW��LT���H��xK���J��xL��XI��    0123456789      basic_string::_M_create %s: __pos (which is %zu) > this->size() (which is %zu)  basic_string::at: __n (which is %zu) >= this->size() (which is %zu) basic_string::erase basic_string::_M_replace_aux basic_string::insert basic_string::replace basic_string::_M_replace basic_string::assign basic_string::append basic_string::copy basic_string::compare     basic_string::_M_construct null not valid basic_string::basic_string string::string basic_string::substr        C POSIX basic_string::erase     %s: __pos (which is %zu) > this->size() �      (which is %zu)  ����h���H���(�����������t���T���4�������%.*Lf %m/%d/%y %H:%M %H:%M:%S   ��� �������������������������������� ��������������� ��0!�� "�����������P"������"��������������������%���%���&���&���'���������%��������������)���(�����������������������������@������j���m��zl��fm��ik��,_��Fb��&a��b��`��    basic_string::_M_create %s: __pos (which is %zu) > this->size() (which is %zu)  basic_string::at: __n (which is %zu) >= this->size() (which is %zu) basic_string::erase basic_string::_M_replace_aux basic_string::insert basic_string::replace basic_string::_M_replace basic_string::assign basic_string::append basic_string::copy basic_string::compare     basic_string::_M_construct null not valid basic_string::basic_string string::string basic_string::substr        std::bad_alloc  std::bad_cast   std::bad_typeid __gnu_cxx::__concurrence_lock_error     __gnu_cxx::__concurrence_unlock_error   std::exception std::bad_exception               0j���j���j���j���      0j��Mk��Mk��Mk��Mk���j��@k���j��0j��            __gnu_cxx::__concurrence_lock_error     __gnu_cxx::__concurrence_unlock_error   __gnu_cxx::__concurrence_broadcast_error        __gnu_cxx::__concurrence_wait_error             pure virtual method called
     deleted virtual method called
  terminate called recursively
   terminate called after throwing an instance of ' '
     terminate called without an active exception
   what():                 rb w+b w r r+ w+ a+ a+b wb ab r+b a u���t��u��u��u���t��u��u��u��\t��u��u���t��lt��u��u���t���t��u��u��|t���t��u��u���t��\t��u��u���t��lt��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u��u���t��u��u��u��|t��u��u��u���t��u��u��u���t��        C       locale::facet::_S_create_c_locale name not valid LC_CTYPE LC_NUMERIC LC_TIME LC_COLLATE LC_MONETARY LC_MESSAGES �����������������������������      ����������      -+xX0123456789abcdef0123456789ABCDEF -+xX0123456789abcdefABCDEF -0123456789 G M T   H S T   A K S T   P �      S T   M S T   C S T   E S T   A S T   N S T   C E T   I S T   E E T   J S T   GMT HST AKST PST MST CST EST AST NST CET IST EET JST      basic_string::replace   %s: __pos (which is %zu) > this->size() (which is %zu)  %m/%d/%y %H:%M:%S  AM PM Sunday Monday Tuesday Wednesday Thursday Friday Saturday Sun Mon Tue Wed Thu Fri Sat January February March April May June July August September October November December Jan Feb Mar Apr Jun Jul Aug Sep Oct Nov Dec % m / % d / % y   % H : % M : % S     A M   P M   S u n d a y   M o n d a y   T u e s d a y   W e d n e s d a y   T h u r s d a y   F r i d a y   S a t u r d a y   S u n   M o n   T u e   W e d   T h u   F r i   S a t   J a n u a r y   F e b r u a r y   M a r c h   A p r i l   M a y   J u n e   J u l y   A u g u s t   S e p t e m b e r   O c t o b e r   N o v e m b e r   D e c e m b e r   J a n   F e b   M a r   A p r   J u n   J u l   A u g   S e p   O c t   N o v   D e c   iostream iostream error Unknown error basic_string::append :    generic system  �      std::bad_array_new_length                       ������������������������������������p���p�������p���p���p���p���p���p���p���p���p���p���p���p�������u���u���u���u���u���u���u���u�������p���p���p���p���p�������p���u�������������������u���u���������������p���p���p�����������������������p�����������p���������������p���p���p���������������p���p���p�������u�������u���u���	���.���.���.���C���	���	��� ��� ���.���.���.���.���.���.���.���.���.���.���.���.���.���.���.���	���.���.���.���.���.���.���.���.���.���.��� ��� ���.���.���	���.���.���.���.������.���.���.���.���	��� ���.���.���.���.���.���.���.���.���.���.���.���.���.���	���	���.���������������	���.���.���.���.���.���.���.���.���(anonymous namespace)   �������������������(������	���	�������������������������������������������������������������������������������������������������������������������������������������������������������������������	�������������������������������������������������������������������������������������������������      st sP cl dt pt qu string literal std auto decltype(auto)    ����������������������������������������������������������������������������L��������������������������������������������������|�����������L�������l������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������o���������������������������������������������������E�������������������������U���=�����������������������������������������o�����������li  ���d���l�������T���\�������"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"�������"���U���"���@���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"���"�������H���Z���Z���(���Z��������������Z���Z���Z���Z���Z���Z���Z���Z�������x���Z���X���8���Z���Z���Z���Z���Z���Z���Z���Z���Z���Z���Z�������Z���Z���Z���Z�������Z���Z���Z���Z���Z���Z���Z���Z���Z���Z���Z���Z���Z�������[abi: :: {default arg# %�      d }:: JArray [] auto: vtable for  VTT for  construction vtable for  -in- typeinfo for  typeinfo name for  typeinfo fn for  non-virtual thunk to  virtual thunk to  covariant return thunk to  java Class for  guard variable for  TLS init function for  TLS wrapper function for  reference temporary #  for  hidden alias for  transaction clone for  non-transaction clone for  _Sat  _Fract _Accum ,  operator operator  ad sZ gs >( ix  :  new  ul ll ull false true java resource  decltype ( ... {parm# this global constructors keyed to  global destructors keyed to  {lambda( )# {unnamed type#  [clone   ����L���L�����������Y�����������)�����,���������������������9�������9�������9�������9���6�������������������������������������������9���9������������ ��� ��y������)���.���)���b���b�����������������������������������d���������������������������)�������i�������i�����������k��������������Y ��������������������w��]��C��1 �� restrict  volatile  const  transaction_safe  noexcept  throw && complex  imagin�      ary  ::*  __vector( �&��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-���)��$*���*���)��$*���*���&���&��$'��d'���(��$+��D(��$)��$-��$-��$-��$-���%��$-���'��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-��$-���,��$-���+��$,�� ( (... ...) _GLOBAL_                          std::allocator allocator std::basic_string basic_string std::string std::basic_string<char, std::char_traits<char>, std::allocator<char> > std::istream     std::basic_istream<char, std::char_traits<char> > basic_istream std::ostream    std::basic_ostream<char, std::char_traits<char> > basic_ostream std::iostream   std::basic_iostream<char, std::char_traits<char> > basic_iostream               t       IaJ            IaJ                            a       �jJ            �jJ            �jJ     	       b       �jJ            �jJ            �jJ            s       �jJ            �jJ     F       �jJ            i       kJ     �             0kJ     1       bkJ            o       pkJ            �kJ     1       �kJ            d       �kJ            �kJ     2       lJ            aN &= aS = aa & an at alignof  az cc const_cast () cm , co ~ dV /= da delete[]  dc dynamic_cast de * dl delete  ds .* . dv / eO ^= eo ^ eq == fL fR fl fr ge >= gt > lS <<= le <= operator""  ls << lt < mI -= mL *= mi - ml mm -- na new[] ne != ng nt ! nw new oR |= oo || or | pL += pl + pm ->* pp ++ ps -> ? rM %= rS >>= rc reinterpret_cast rm % rs >> sizeof... sc static_cast sizeof  sz tr throw tw throw     �mJ     �mJ           �mJ     �mJ           �mJ     iJ           �fJ     �mJ           �mJ     �mJ           �mJ     �mJ           �mJ     �mJ           �mJ     �mJ     
      .aJ     �mJ           �mJ     �mJ           �mJ     �mJ           �mJ     �mJ           �mJ     �mJ     	      �mJ     �mJ           nJ     nJ           nJ     nJ           nJ     nJ           1aJ     nJ            nJ     #nJ           �      %nJ     (nJ           +nJ     .nJ           0nJ     3nJ           6nJ     gJ           9nJ     gJ           <nJ     gJ           ?nJ     gJ           BnJ     EnJ           �fJ     eJ           HnJ     KnJ           �fJ     -eJ           MnJ     PnJ           TnJ     WnJ           TcJ     ZnJ           fnJ     inJ           lnJ     onJ           qnJ     tnJ           wnJ     znJ           }nJ     �nJ           �nJ     nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           4aJ     �nJ           7aJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ           �nJ     �nJ            oJ     oJ           +aJ     oJ     	      �fJ     �      oJ     	      oJ     oJ           (aJ     oJ           'oJ     oJ           *oJ     -oJ            3oJ     6oJ                                   signed char bool boolean char byte double long double float __float128 unsigned char int unsigned int unsigned long unsigned long __int128 unsigned __int128 short unsigned short void wchar_t long long unsigned long long decimal32 decimal64 decimal128 half char16_t char32_t decltype(nullptr)                             �uJ            �uJ            �uJ            �uJ           �uJ            �uJ            �uJ            �uJ           �uJ            �uJ           �uJ            �uJ           �uJ     
       �uJ     
      �uJ            �uJ            �uJ            �uJ           �uJ            vJ                                           vJ            vJ           vJ            vJ           "vJ            "vJ            +vJ            +vJ                                                                    �                                              =vJ            =vJ            CvJ            CvJ                                            RvJ            RvJ        	   WvJ            �uJ            _vJ     	       vJ           ivJ            ivJ           gJ            gJ            |vJ     	       |vJ     	       �vJ     	       �vJ     	       �vJ     
       �vJ     
       �vJ            �vJ           �vJ            �vJ            �vJ            �vJ            �vJ            �vJ            `�L     ��L                     ��@                               M      M     �L     @M                                     Argument domain error (DOMAIN) Argument singularity (SIGN)      Overflow range error (OVERFLOW) Partial loss of significance (PLOSS)    Total loss of significance (TLOSS)      The result is too small to be represented (UNDERFLOW) Unknown error     _matherr(): %s in %s(%g, %g)  (retval=%g)
  �5��5���5���5���5���5���5��Mingw-w64 runtime failure:
     Address %p has n�      o image-section   VirtualQuery failed for %d bytes at address %p          VirtualProtect failed with code 0x%x    Unknown pseudo relocation protocol version %d.
         Unknown pseudo relocation bit size %d.
               .pdata          �M���M���M��N���M��pM���M��    �N��pN��`N��@N���N��pN��        INF INITY NAN                   Lɚ� �R`�%uM��]=�];���Zeu��uv�HMe�Ƒ����F�ݍ�����~�QCo�ߌ��G���A�<զ��Ix��@ �p+��ŝi@     ���4@        ��@        @�@         �@         �@             ��?                    alnum alpha cntrl digit graph lower print punct space upper xdigit                               J           J           J             J            J           J            $J     W      *J            0J            6J            <J     �                                                        	               	      
                                                !      5      A      C      P      R      S      W      �      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �               ����                nf inity an f��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��$g��$g��$g��$g��$g��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��$g��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��Dg��tf��Dg��g��                                         
                              !   #   &   (   *   -   /   1   4             �?               @      �?  �����AV瞯�<       �        (null) NaN Inf  ( n u l l )     p���������������������������������������@���s�������í��#�������б�������������������������������������������������������������������������Ұ���������@���s��������������������������������������������� �������������������d������������������������������������������0�������@������������������Я������s���`��� ���d��������������� ���Я��d�����������d�������Я��    Infinity NaN 0  ���$���$���b���5���          �?�      aCoc���?��`�(��?�y�PD�?�}�-�<2ZGUD�?      �?      $@      @      @      @       �              �?        ABCDEF abcdef 0123456789                              }                             �?      $@      Y@     @�@     ��@     j�@    ��.A    �cA    �חA    e��A    _�B   �vH7B   ��mB  @�0�B  �ļ�B  4&�kC ��7y�AC �؅W4vC �Ngm��C =�`�X�C@��x�DP����KD��M���D        ��ؗ�Ҝ<3���#�I9=��D��2�����[%Co�d(�
                         ��7y�ACn����F��?�O8M20�Hw�Z<�s�Ou                        C%p %d %s
 C%p %d V=%0X w=%ld %s
               %p not found?!?!
       Error cleaning up spin_keys for thread                                                                      once %p is %d
 T%p %d %s
 T%p %d V=%0X H=%p %s
             ../../src/mingw-w64/mingw-w64-libraries/winpthreads/src/rwlock.c        (((rwlock_t *)*rwl)->valid == LIFE_RWLOCK) && (((rwlock_t *)*rwl)->busy > 0)    Assertion failed: (%s), file %s, line %d
 RWL%p %d %s
  RWL%p %d V=%0X B=%d r=%ld w=%ld L=%p %s
        PJ     �              �J             �J             �J             �'J             @(J             �(J              )J             `)J             �)J              *J             �*J             �+J             `,J              -J             �-J             �.J             �.J             ��F             @�J              /J             /J              /J             0/J             @/J             P/J             `/J             дF             �F             ��F             ��F             `�F             �G             ��G             �#H             �GH             �SH              1J             �1J             ��H              2J             02J             @2J             �J              �J             �2J             �2J             �2J             �2J             �2J             �2J             �2J             �2J              3J             3J              3J             03J             @3J             P3J             `3J             p3J             �3J             �3J             �3J             �      �3J             �3J             �3J             �3J             �3J              4J             4J              4J             04J             0[I             @4J             P4J             `4J             p4J             �4J             �4J             �4J             �4J             �4J             �4J              �I             �4J             �4J              5J             5J              5J             @6J             `7J             �8J             �I             �9J             �:J             �;J              =J             �J             0�J             ��J              �J             p�J             ��J             P�J             ��J              �J             ��J             0�J             ��J             ��J             @ K             p K             � K             � K             �K             0K             �K             �K              K             �K              K             �K             �K             �K              K             PK             �K     �              K             �K             	K             `	K             �	K             �K              K             �K             K             �K             �K              K             0K             `K             �K             �K             �K             �K             �K             �K             K             0K             �K             �K             �K             @K             �K             �K              K              K             `K             �K              K             �K              K             `K             0K             �K             �K               K             p K             � K             � K              !K              !K             p!K             �!K             �!K              "K              J              %K              %K             ��J              {J             @�L               @             ��L             ��L             ��L             �L             `�L             0�L             8�L             �      ��J             `�J              M             M             M             0M             0J             P�L             �@             ��@              �L             0�L             `�L             �L             �L             �L             ?                          YXJ     bXJ     mXJ     uXJ     �XJ     �XJ                     �������                        ��������        �������?                        ��������                                                                                                                @                                                                                                                                                       ��              ﻿             ��                                                                                           ��J             �4J      3J     �3J     �2J     �4J     @3J     �4J     `3J      5J     �3J     /J     �2J      /J     �2J     `4J      3J     �4J     03J     �3J     �      �2J     �4J     P3J     �4J     p3J     5J     �3J     0/J     �2J     @/J     �2J     p4J     3J                                     ?                                                              P/J     @3J     �4J     `/J     P3J     �4J                      2J     �3J     02J     �3J     �3J     �3J                     �2J     �2J                      4J      4J      3J     4J     04J     03J                      3J     3J                     `3J     �3J     �2J     �2J     p3J     �3J     �2J     �2J                                     ��J      �J      �J     ��J     ��J     `�J                                    C                                                                                                                                          ��������        ��������                                                                                                   �                                                                                                          �                                    @                                                             �                                                                                                                                                                                       J                                              @                                             �J                     �����������������J                                     �J                     ���������������� �J                     �               ��J                     �       ����������J                     (�������(���������J                             �               �J                     (�������(��������J                     �                �J                     8�������8������� �J                     �               ��J                     (�������(���������J                     �               p�J                     �       ��������p�J                     (�������(�������p�J                     �              �               еJ                     8�������8�������еJ                     �               �J                     0�������0��������J                     �               ��J                     0�������0���������J                                    ��J                     ������������������J                                    еJ                     ����������������еJ                     �                �J                     8�������8������� �J                     �               еJ                     8�������8�������еJ                      �J     ��J     ��J     ��J     ��J              �J      �J     ��J     `�J     �J             ��J     ��J     �J             ��J     ��J     ��J             ��J      �J     ��J             ��J     `�J     ��J             ��J     ��J      �J             ��J     ��J     @�J             ��J      �J     ��J             ��J     `�J     ��J             ��J     ��J     �J             ��J     ��J     �J             ��J      �J     �J             �      ��J     `�J     �J             ��J     ��J            @�J            ЬJ                   ��J     ��J            p�J            ЬJ                   ��J      �J            `�J            ЬJ                   ��J     `�J            ��J            ЬJ                   ��J     ��J            0�J            ЬJ                    ��J     ��J            ��J            ЬJ                    ��J      �J            p�J            ЬJ                    ��J     `�J            �J            ЬJ                    ��J     ��J            ��J            ЬJ                   ��J     ��J            0�J            ЬJ                   ��J      �J            пJ            ЬJ                   ��J     `�J            P�J            ЬJ                   ��J     ��J            �J            ЬJ                   ��J     ��J            p�J            ЬJ                   ��J      �J            0�J            ЬJ                   ��J     `�J            �      ��J            ЬJ                   ��J     ��J             �J            ЬJ                   ��J     ��J            �J            ЬJ                   ��J      �J            @�J            ЬJ                   ��J     `�J            �J            ЬJ                   ��J     ��J            `�J            ЬJ                   ��J     ��J            0�J            ЬJ                   ��J      �J            ��J            ЬJ                   ��J     `�J            P�J            ЬJ                   ��J     ��J            ��J            ЬJ                   ��J     ��J            �J            ЬJ                   ��J      �J            вJ            ЬJ                   ��J     `�J            0�J            ЬJ                   ��J     ��J            �J            ЬJ                   ��J     ��J            p�J            ЬJ                   ��J      �J            P�J            ЬJ                   ��J     `�J     �             ��J            ЬJ                    �J     ��J      �J     ��J      �J     ��J     ��J      �J            �J            ��J                    ��J      �J            �J            ��J                    ��J     @�J            �J            ��J                    ��J     `�J            �J            ��J                    ��J     ��J     p�J             ��J     ��J     ��J             ��J     ��J     ��J             ��J      �J     �J             ��J     @�J     0�J             ��J     ��J     P�J             ��J     ��J     p�J             ��J      �J     ��J             ��J     ��J     �J             ��J     ��J     0�J             ��J      �J     p�J             ��J     @�J     ��J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J            �J             �J                    ��J     ��J            �J             �J                    ��J      �J     �J             ��J      �J     �J             ��J     @�J            �      �J            ��J                    ��J     ��J            �J            ��J                    ��J      �J     �J             ��J     `�J     �J             ��J     ��J     �J             ��J      �J     �J             ��J     ��J     ��J             ��J     ��J     �J             ��J     ��J           �J             �J                   ��J     ��J            ��J     �������        ��J     ��J            ��J     �������        ��J     ��J     �J              �J      �J      �J     �J     ��J      �J            �J            ��J                    ��J     @�J            �J            ��J                    ��J     `�J            �J            ��J                    ��J     ��J            �J            ��J                    ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J              �J      �J     ��J      �J     `�J             ��J     @�J     ��J             ��J     `�J     гJ             �      ��J     ��J     гJ             ��J     ��J     гJ             ��J     ��J     �J             �K     ��J     p�J             ��J      �J     �J             ��J      �J     ��J             ��J     `�J     ��J             ��J     ��J     ��J             ��J     ��J     p�J             ��J      �J            ��J     �������        ��J     `�J            ��J     �������         �J     ��J     ��J     ��J     �J             ��J     ��J     �J             ��J      �J     ��J             ��J     `�J           ��J            еJ                   ��J     ��J      �J             ��J     ��J     еJ             ��J      �J      �J             ��J     @�J      �J             ��J     `�J     @�J             ��J     ��J     `�J             ��J     ��J     �J              �J     ��J      �J      �J     ��J     @�J     0�J             ��J     `�J     p�J             ��J     ��J     ��J             ��J     ��J     пJ             ��J     ��J     �J             ��J      �J     0�J             ��J     �      ��J     p�J             ��J     ��J     ��J             ��J     @�J     �J             ��J     `�J     �J             ��J     ��J     �J             ��J     ��J     гJ             ��J     ��J     �J             ��J     ��J     �J             ��J      �J     ��J             ��J      �J     вJ             ��J     @�J     �J             ��J     `�J     P�J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J             ��J      �J     ��J             ��J      �J     �J             ��J     @�J      �J             ��J     `�J             �J                     ��J     ��J     ��J             ��J     ��J     �J             ��J     ��J      �J             ��J     ��J     ��J             ��J      �J            �J            p�J                    ��J      �J            �J            p�J                    ��J     @�J            �J            �J                    ��J     ��J            �J            �J     �                     ��J     ��J            �J            �J                    ��J      �J            �J            �J                    ��J     @�J     ��J             ��J     ��J     �J             ��J     ��J      �J             ��J      �J            �J            p�J                    ��J     �J     ��J             ��J      �J      �J             ��J     @�J     @�J             ��J     `�J     ��J             ��J     p�J     ��J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J             ��J     ��J     �J             ��J      �J     �J             ��J     `�J     �J             ��J     ��J     �J              �J     ��J     ��J     ��J            �J             �J                    ��J     ��J            �J             �J                    ��J     ��J     �J             ��J     ��J     �J             ��J      �J            �J            ��J                    ��J     @�J            �J            ��J            �              ��J     ��J     �J             ��J     ��J     �J             ��J      �J     �J             ��J      �J      �J             ��J     `�J      �J              �J     ��J     ��J     ��J     �J             ��J      �J     �J             ��J     @�J     �J             ��J     ��J     �J              �J     ��J      �J     ��J     N10__cxxabiv115__forced_unwindE N10__cxxabiv117__class_type_infoE                               N10__cxxabiv119__foreign_exceptionE                             N10__cxxabiv120__si_class_type_infoE                            N10__cxxabiv121__vmi_class_type_infoE                           *N12_GLOBAL__N_117io_error_categoryE                            *N12_GLOBAL__N_121system_error_categoryE                        *N12_GLOBAL__N_122generic_error_categoryE                       N9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE                N9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE                N9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE           �      N9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE           N9__gnu_cxx24__concurrence_lock_errorE                          N9__gnu_cxx24__concurrence_wait_errorE                          N9__gnu_cxx26__concurrence_unlock_errorE                        N9__gnu_cxx29__concurrence_broadcast_errorE                     *NSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE             *NSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE             *NSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE             *NSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE             *NSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE            *NSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE            *NSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE    �              *NSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE            *NSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE            *NSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE            *NSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE            *NSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE           *NSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE           *NSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE           *NSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE           *NSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE           *NSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE           *NSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE           *NSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE           *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_sh�      imIcLb1EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE      *NSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE      NSt3_V214error_categoryE        NSt6locale5facet6__shimE        NSt6locale5facetE               NSt7__cxx1110moneypunctIcLb0EEE NSt7__cxx1110moneypunctIcLb1EEE NSt7__cxx1110moneypunctIwLb0EEE NSt7__cxx1110moneypunctIwLb1EEE NSt7__cxx1114collate_bynameIcEE NSt7__cxx1114collate_bynameIwEE NSt7__cxx1115messages_bynameIcEE                                NSt7__cxx1115messages_bynameIwEE                                NSt7__cxx1115numpunct_bynameIcEE                                NSt7__cxx1115numpunct_bynameIwEE                                NSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE                    NSt7__cxx1115time_get_bynameIwSt19istrea�      mbuf_iteratorIwSt11char_traitsIwEEEE                    NSt7__cxx1117moneypunct_bynameIcLb0EEE                          NSt7__cxx1117moneypunct_bynameIcLb1EEE                          NSt7__cxx1117moneypunct_bynameIwLb0EEE                          NSt7__cxx1117moneypunct_bynameIwLb1EEE                          NSt7__cxx117collateIcEE         NSt7__cxx117collateIwEE         NSt7__cxx118messagesIcEE        NSt7__cxx118messagesIwEE        NSt7__cxx118numpunctIcEE        NSt7__cxx118numpunctIwEE        NSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE                            NSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE                            NSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE                           NSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE                           NSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE                           NSt7__cxx119money_putIwSt19ostre�      ambuf_iteratorIwSt11char_traitsIwEEEE                           NSt8ios_base7failureB5cxx11E    NSt8ios_base7failureE           Sd              Si              So              St10bad_typeid  St10ctype_base  St10money_base  St10moneypunctIcLb0EE           St10moneypunctIcLb1EE           St10moneypunctIwLb0EE           St10moneypunctIwLb1EE           St11__timepunctIcE              St11__timepunctIwE              St11logic_error St11range_error St12codecvt_base                St12ctype_bynameIcE             St12ctype_bynameIwE             St12domain_error                St12length_error                St12out_of_range                St12system_error                St13__ios_failure               St13bad_exception               St13basic_filebufIcSt11char_traitsIcEE                          St13basic_filebufIwSt11char_traitsIwEE                          St13basic_fstreamIcSt11char_traitsIcEE                          St13basic_fstreamIwSt11char_traitsIwEE                          St13basic_istreamIwSt11c�      har_traitsIwEE                          St13basic_ostreamIwSt11char_traitsIwEE                          St13messages_base               St13runtime_error               St14basic_ifstreamIcSt11char_traitsIcEE                         St14basic_ifstreamIwSt11char_traitsIwEE                         St14basic_iostreamIwSt11char_traitsIwEE                         St14basic_ofstreamIcSt11char_traitsIcEE                         St14basic_ofstreamIwSt11char_traitsIwEE                         St14codecvt_bynameIcciE         St14codecvt_bynameIwciE         St14collate_bynameIcE           St14collate_bynameIwE           St14overflow_error              St15basic_streambufIcSt11char_traitsIcEE                        St15basic_streambufIwSt11char_traitsIwEE                        St15messages_bynameIcE          St15messages_bynameIwE          St15numpunct_bynameIcE          St15numpunct_bynameIwE          St15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE                              St15time_get_byn�      ameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE                              St15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE                              St15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE                              St15underflow_error             St16__numpunct_cacheIcE         St16__numpunct_cacheIwE         St16invalid_argument            St17__timepunct_cacheIcE        St17__timepunct_cacheIwE        St17moneypunct_bynameIcLb0EE    St17moneypunct_bynameIcLb1EE    St17moneypunct_bynameIwLb0EE    St17moneypunct_bynameIwLb1EE    St18__moneypunct_cacheIcLb0EE   St18__moneypunct_cacheIcLb1EE   St18__moneypunct_cacheIwLb0EE   St18__moneypunct_cacheIwLb1EE   St19__codecvt_utf8_baseIDiE     St19__codecvt_utf8_baseIDsE     St19__codecvt_utf8_baseIwE      St19__iosfail_type_info         St20__codecvt_utf16_baseIDiE    St20__codecvt_utf16_baseIDsE    St20__codecvt_utf16_baseIwE     St20bad_array_new_length        St21__ctype_abstract_baseIcE    St21__ct�      ype_abstract_baseIwE    St23__codecvt_abstract_baseIDiciE                               St23__codecvt_abstract_baseIDsciE                               St23__codecvt_abstract_baseIcciE                                St23__codecvt_abstract_baseIwciE                                St25__codecvt_utf8_utf16_baseIDiE                               St25__codecvt_utf8_utf16_baseIDsE                               St25__codecvt_utf8_utf16_baseIwE                                St5ctypeIcE     St5ctypeIwE     St7codecvtIDiciE                St7codecvtIDsciE                St7codecvtIcciE St7codecvtIwciE St7collateIcE   St7collateIwE   St7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE       St7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE       St7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE       St7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE       St8bad_cast     St8ios_base     St8messagesIcE  St8messagesIwE  St8numpunctIcE  St8numpunctIwE  St8time_getIcSt19istreambuf_iter�      atorIcSt11char_traitsIcEEE      St8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE      St8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE      St8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE      St9bad_alloc                    St9basic_iosIcSt11char_traitsIcEE                               St9basic_iosIwSt11char_traitsIwEE                               St9exception                    St9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE     St9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE     St9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE     St9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE     St9time_base    St9type_info    xK     8�J     `�J     ��J     ��J     �K     �K             �K      K     HK     pK     (K     ؞J     X�J     ��J     ��J     ПJ     (�J      �J     xK     PK     �K     H�J     ��J      �J     ȠJ     �J     ��J     p�J     �K     �K     (	K     P	K     x	K     �	K     �	K     �J     @�J     �       
K     H
K     h�J     ��J     p
K     �
K     ��J     �J     �J     0�J     �
K     �
K             K     X�J     ��J     @K     hK     ��J     ТJ     �K             �J                     `J                     �J     0�A      �A     p�E     p�E      �A     ��A     P�A     ��A     `�A                     �J                     `J                      �J     ��A     `�A     p�E     p�E      �A     ��A     p�A     ��A     ��A                     @�J     ��A     ��A     p�E     p�E      �A     ��A     0�A     P�A     ��A                     `�J     @�A     �A     ��A     @`B     ��A     �aB     PaB     0aB             ��J     `�A     P�A     @�A     @`B     `�A     �aB     PaB     0aB             ��J     ��A     ��A     P�A     @`B     `�A     �aB     PaB     0aB             ��J     ��A     ��A     �!G     �#G     @(G     *G     ` G     �-G     $G     �.G     0&H     �,G     P&G     �*G             �J     ��A     ��A     �DG     GG     �KG     PMG     �CG     PQG     pGG      RG     �       0H      PG     �IG      NG              �J     ��A     `�A     p%H     �&H     P�A     ��A     ��A     P+H     ��A     ��A     ��A     ��A     0�A     P�A              �J     `�A     0�A     p/H     �0H     ��A     P�A     ��A     @5H     �A     `�A     ��A      �A     ��A     ��A             @�J     ��A     ��A     ��A                     `�J     0�A      �A     ��A                     ��J     p�A     @�A     ��A                     ��J     ��A     ��A     ��A                     ��J     �F     p�F      )B     `)B     `�C                      �J     `�F     ��F     0)B     �)B      �B                     @�J     P�F     ��F     �*B     �*B     P�C                     ��J     ��F      �F     �*B     �+B     `�B                     ��J     p�F     ��F     �-B     �,B      .B                      �J     ��F     0�F     �-B      ,B     .B                     @�J     P�F     ��F     �/B     �.B      0B                     ��J     ��F     �F     �/B      .B     0B                     ��J     P�F     �      ��F     �E     �E     �E     E     @E                      �J     ��F      �F     `�B     p�B     �B     `�B     ��B                     @�J     p�F     ��F     � E     � E     �E      E     @ E                     ��J     ��F      �F      �B     0�B     нB      �B     p�B                     ��J     ��F     ��F     �2B      1B      0B     �2B     �3B     �1B              �J     ��F     @�F     �2B     p1B     �0B     P3B     04B     P2B     `�B                     @�J     ��F     �F     @7B     �5B     �4B     `7B     @8B     `6B             ��J     ��F     `�F     P7B     �5B     5B     �7B     �8B     �6B     P2C                     ��J     ��F     0�F      =B     @;B              �J     �F     ��F     �=B      9B             @�J     ��F     P�F     �BB      AB             ��J     0�F     ��F     �CB     �>B             ��J     �F     p�F     �FB     �EB              �J     P�F     ��F     @GB     �DB             @�J     0�F     ��F     �IB     �HB             ��J     p�F     ��F     �      0JB     �GB             ��J     ��F     ��F     �B      B     �B     pB     �B     �B     �B     �B     �B                      �J     ��F      �F     ��B     ��B     ��B     ��B     P�B      �B     ��B     p�B     `�B                     @�J     0�F     P�F     �B     `B     0B     �B     0B      B     �B     �B     �B                     ��J     ��F     ��F     0�B     ��B     ��B     ЊB     ��B     @�B      �B     ��B     ��B                     ��J     ��F     ��F     0B     �B     pB     �B     pB     @B      B     B      B                      �J     0�F     `�F     p�B      �B     0�B     �B     ЏB     ��B     `�B     ��B     ��B                     @�J     p�F     ��F     pB     �B     �B     0B     �B     �B     `B     PB     @B                     ��J     ��F      �F     ��B     `�B     p�B     P�B     �B     ��B     ��B     0�B      �B                     ��J                     `J     @`B     `J     �aB     PaB     0aB             �J     ��H     �      ��H             �J     �H     ��H     ��B     ��B     ��B     ��B     P�B      �B     ��B     p�B     `�B                     0�J     ��H     p�H     0�B     ��B     ��B     ЊB     ��B     @�B      �B     ��B     ��B                     p�J     p�H     @�H     p�B      �B     0�B     �B     ЏB     ��B     `�B     ��B     ��B                     ��J     @�H     �H     ��B     `�B     p�B     P�B     �B     ��B     ��B     0�B      �B                     �J     0 I       I     ��B     �B      �B                     �J     @$I     $I     ��B     �B     `�B                     0�J     P&I      &I     ��B     ��B     йB                     P�J     `(I     0(I     �B     ��B      �B                     p�J     p,I     @,I     `�B     p�B     �B     `�B     ��B                     ��J     @0I     0I      �B     0�B     нB      �B     p�B                     ��J     1I     �0I     `�B      �B     ��B     �B     0�B     @�B     `�B                     ЮJ     �1I     �1I     0C     `�B     �      ��B     �C     C     ��B     P2C                     �J     �5I     �5I     ��B     ��B     ��B     ��B     P�B      �B     ��B     p�B     `�B                     �J     �9I     P9I     0�B     ��B     ��B     ЊB     ��B     @�B      �B     ��B     ��B                     0�J     P=I      =I     p�B      �B     0�B     �B     ЏB     ��B     `�B     ��B     ��B                     P�J      AI     �@I     ��B     `�B     p�B     P�B     �B     ��B     ��B     0�B      �B                     p�J     �BI     `BI     ��B     �B      �B                     ��J     @DI     DI     ��B     �B     `�B                     ��J     FI     �EI     ��B     ��B     йB                     �J     �GI     �GI     �B     ��B      �B                     0�J     �KI     PKI     `�B     p�B     �B     `�B     ��B                     P�J     �NI     �NI      �B     0�B     нB      �B     p�B                     p�J     �OI     �OI     `�B      �B     ��B     �B     0�B     @�B     `�B                     �      ��J     @PI     PI     0C     `�B     ��B     �C     C     ��B     P2C                     �J     �PI     �PI     XC     0VC             �J     `QI     0QI     p{C     �yC             0�J     �QI     �QI     ~C     �}C             P�J     �RI     PRI     @�C     ��C             p�J     tI     �sI     pE                     ��J     �tI     ptI     `E                            ��J     �F     0F            ����������J     ��I     ��I     ������������������J     ��I     P�I                            �J     �JF     �JF     �����������������J     @�I     ��I                     �J     �nF     `nF     ���������������� �J     ��I     p�I             P�J     ��F     `�F     �B                     ��J      �F     �F     �B      B     �B     pB     �B     �B     �B     �B     �B                     вJ     ��F     ��F     �B     `B     0B     �B     0B      B     �B     �B     �B                     �J     ��F     ��F     0B     �B     pB     �B     pB     @B     �       B     B      B                     P�J     ��F     P�F     pB     �B     �B     0B     �B     �B     `B     PB     @B                     ��J     ��F     `�F             ��J     �F     вF             гJ     дF     ��F     �(B                     �J     �F     ��F     @KB                      �J     ��F     ��F     �bB     @bB      bB     �aB      eB     �dB     0eB     eB             @�J     ��F     ��F     phB     �gB     @eB     PfB     @fB     �eB     �eB     �eB     iB     �hB      jB      iB             `�J     ��F     ��F     �(B                     ��J     ��F     p�F     �(B                     ��J     `�F     0�F     �(B                     ��J     ��F     p�F     @KB                     �J     0G     �G     pE                      �J     �G     pG     �JB                      �J     �9G     �9G     �!G     �#G     @(G     *G     ` G     �-G     $G     �.G     0&H     �,G     P&G     �*G             @�J     p]G      ]G     �DG     GG     �KG     PMG     �CG     �      PQG     pGG      RG      0H      PG     �IG      NG     �               `�J     �lG     @lG     �       ��������`�J     ��I      �I     (�������(�������`�J     ��I     ��I             �               ��J     �|G     �{G     �       ����������J      �I     p�I     (�������(���������J     ��I     @�I                            ��J      �G     ��G     ������������������J     ��I     ��I                    еJ     p�G     0�G     ����������������еJ     `�I      �I             �J     ��G     p�G     @KB             �               0�J     ��G     P�G     0�������0�������0�J     0�I     ��I     �               P�J     ��G     P�G     0�������0�������P�J     `�I     ��I                    p�J      �G     ��G            ��������p�J     �I     ��I     ����������������p�J     P�I     ��I             �               ��J     �H     0H     8�������8���������J      �I     ��I     �               жJ      H     pH     8�������8�������жJ     @�I     ��I             �J     �H     pH     ��C     `�C     �      ��C     p�C     ��C     ��C     p�C                     �J     �H     �H      �C     `�C     0�C     ��C      �C     P�C     �C                     0�J     �H     PH      �C     p�C     `�C                     P�J     �"H     `"H     �C     0�C     P�C                     p�J     �#H     p#H     @KB                     ��J      -H     �,H     p%H     �&H     �)H      *H     P%H     P+H     0(H     �+H     0&H     +H     )H     �*H             ��J     7H     �6H     p/H     �0H     �3H     �3H     P/H     @5H      2H     �5H      0H      5H      3H     �4H             ��J     P9H      9H     �E     pE     �E                     зJ     `;H     0;H     �E     �E     �E                     �J     p?H     @?H     �E     �E     �E     E     @E                     �J     @CH     CH     � E     � E     �E      E     @ E                     0�J     DH     �CH     �&E     P#E     "E     `*E     �/E     �$E             P�J     �DH     �DH     �\E     �XE     0WE     �_E     `eE     �      PZE             p�J     �EH     �EH      �E                     ��J      GH     �FH     ��E                     ��J     �GH     �GH     @KB                     иJ     �LH     �LH             �J     `RH     0RH             �J     �SH     �SH     �(B                     0�J     XH     �WH             P�J     `\H     0\H             p�J     0`H      `H     �B      B     �B     pB     �B     �B     �B     �B     �B                     ��J      dH     �cH     �B     `B     0B     �B     0B      B     �B     �B     �B                     ��J     �gH     �gH     0B     �B     pB     �B     pB     @B      B     B      B                     йJ     �kH     pkH     pB     �B     �B     0B     �B     �B     `B     PB     @B                     �J     �qH     �qH             �J     �xH     pxH             0�J     �H     �H             P�J     @�H     �H             p�J     0�H      �H     `MB      �C     �LB     0�C     P�C      NB     �LB                     ��J     �      p�H     @�H     0OB      �C     �NB     0�C     P�C     �OB     �NB                     ��J     ��H     ��H     �PB      �C      PB     0�C     P�C      QB     �OB                     кJ     ��H     ��H     p�E     p�E      �A     0QB     p�A     ��A     ��A                      �J     0�H      �H     �UB      �C     PTB     0�C     P�C     �VB     0TB                      �J     p�H     @�H     �WB      �C     PWB     0�C     P�C     PXB     0WB                     @�J     ��H     ��H     0YB      �C     �XB     0�C     P�C     �YB     �XB                     `�J     ��H     ��H     �YB                     ��J                     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J             ��J                     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J     `J              �J                     `J     `J     `J     `J     `J     `J     `J                     @�J                     `J     `J     `J     �      `J     `J     `J     `J                     ��J                     `J     `J     `J     `J     `J     `J     `J                     ��J                     `J     `J     `J     `J     `J     `J     `J                      �J     0�H      �H     @[B      �C      ZB     0�C     P�C     P\B      ZB                      �J     p�H     @�H      ]B      �C     �\B     0�C     P�C     �]B     �\B                     @�J     ��H     ��H      _B      �C     �]B     0�C     P�C     `B     �]B                     `�J     ��H     ��H     �bB     @bB      bB     �aB      eB     �dB     0eB     eB             ��J     ��H     p�H     phB     �gB     @eB     PfB     @fB     �eB     �eB     �eB     iB     �hB      jB      iB             ��J     �RI     �RI      �C      �C     ��C     0�C     P�C     ��C     @�C                     �J     SI     �RI     ЦC      �C     `�C     0�C     P�C     0�C     @�C                      �J     �SI     �SI     ��C     `�C     ��C     p�C     ��C     ��C     �      p�C                      �J      UI     �TI      �C     `�C     0�C     ��C      �C     P�C     �C                     @�J     �VI     �VI      �C     p�C     `�C                     `�J     `XI     0XI     �C     0�C     P�C                     ��J     0YI      YI     �>D     pID     0JD     ID     �ID     �JD     �JD     �GD     �CD     �ED     �=D                     ��J     �YI     �YI     ��D     ��D     P�D     0�D     ��D     ��D     �D     �D     ��D     ��D      �D                     ��J     PZI      ZI     @�D     �E      E     @E     �E     E     `E     ��D             �J     �ZI     �ZI     �E     PE     �E     �E     E     �E     �E     `E              �J     0[I      [I     PE                      �J     �uI     puI             0�J     `wI     0wI     �E     pE     �E                     p�J     0yI      yI     �E     �E     �E                     ��J     �|I     �|I     �E     �E     �E     E     @E                     пJ     @�I     �I     � E     �      � E     �E      E     @ E                     �J      �I     ЀI     �&E     P#E     "E     `*E     �/E     �$E             0�J     ��I     `�I     �\E     �XE     0WE     �_E     `eE     PZE             p�J      �I     ��I      �E                     ��J     ��I     ��I     ��E                     ��J      �I     ЂI     ��E                     ��J     @�I     �I             ��J      �I     �I             �J     P�I     @�I     P�E                      �J     ЕI     ��I      �E     �E             @�J     `�I     0�I     ��E     ��E             `�J     �I     ��I     ��E     @�E             ��J     ��I     P�I     ��E     0�E             ��J     ��I     ��I     p�E     p�E     P�E     `�E                                                     `@@@@@@@@@@@@@@@X X X X X X X X X X @@@@@@@U U U U U U E E E E E E E E E E E E E E E E E E E E @@@@@@V V V V V V F F F F F F F F F F F F F F F F F F F F @@@@                                 �                                                                                                                                                                                                                                      GCC: (x86_64-posix-seh-rev0, Built by MinGW-W64 project) 8.1.0  GCC: (x86_64-posix-seh-rev0, Built by MinGW-W64 project) 8.1.0                                                                                                                                                                                                                                                                        �   !  � 0  y  � �  �  � �  �  (� �    H�   )  h� 0  <  p� @  A  t� P  �  x� �  �  �� �  �  �� �    ��   +  �� +  g  �� g  �  �� �    ��    o  �� p  �  �� �  y  �� �  7  �� @  �  ȹ �  �  й �  H  ع P  �  � �    �     ��    �   � �  �  � �  R  � `  �  � �  �  � �  >    � @   	!  ,� �      !  �"  <� �"  @)  D� @)  �)  X� �)  +  h� +  3+  x� @+  �0  |� �0  �:  �� �:  �<  �� �<  d=  �� p=  �?  �� �?  @  к  @  �@  ܺ �@  �D  �  E  �K  �� �K  
�   � �  ��  � ��  ��  $� ��  ��  8� ��  ��  H�  �  ��  \� ��  9�  p� @�  A�  �� P�  צ  �� �  �  �� �  e�  �� p�  ��  л ��  խ  x� �  F�  �� P�  o�  �� p�  w�  �� ��  ��  �� ��  f�  �� p�  h�  �� p�  ��  �� ��  �  ��  �  #�  ̼ 0�  q�  м ��  ��  ؼ ��  ��  ܼ ��  ��  �� ��  ��  �� ��  ��  �� ��  ��  � ��  K�  � P�  �  4� �  ܹ  <� �  ǻ  L� л  :�  T� @�  ��  d� ��  `�  t� `�  :�  |� @�  ^�  �� `�  r�  �� ��  ľ  �� о  ]�  �� `�  Կ  �� �  �  ��  �  ��  �� ��  ��  �� ��  a�  �� p�  �  Ľ `�  ��  ̽ ��  ��  Խ ��  ��  ܽ  �  �  � �  �  �  �  +�  � 0�  5�  � @�  I�  �� P�  _�  �� `�  ��  �� ��  ��  � ��  ��  � ��  ��  � ��  �   � �  ��  (� ��  ��  8� ��  �  @� �  %�  D� 0�  ��  H� ��  ��  `� ��  �  l� �  ��  t� ��  
�  �� �  ��  �      ��  �  ��  �� ��   �  ��  �  �  �� ��  ��  �� ��  ��  �� ��  8�  о @�  t�  � ��  ��  �� ��  O�  � P�  ��  � ��  ��  � ��  �  0� �  p�  8� p�  u�  D� ��  �  H� �  ��  T� ��  ��  `�  �  ��  x� ��  R�  �� `�  ��  �� ��  ��  �� ��  ��  ��  �  ��  �� ��  4�  �� @�  l�  ̿ p�  ��  п  �  J ؿ P � �� � P � P 2  � @  (�   V ,� ` � 0� � 
 4�  
 5 L� @ y `� � � d� � � p� � � t� � � |� � O �� P � ��   � �� � D �� P [ �� ` ) �� 0 w �� �  ��    ��   � �� � �  � �  n# � p# L$ ,� P$ �$ 8�  % �& D� �& �) P�  * �. h�  / 8 |� 8 @8 �� @8 �8 �� �8 �8 �� �8 �: �� �: P ��  P /Y �� 0Y #Z �� 0Z sZ � �Z [ �  [ �^ � �^ �_ (� �_ �_ 4� �_ �` <� �` Ca H� Pa �a P�  b &b `� 0b Qc h� `c �d |� �d �e �� �e f ��  f �g �� �g �h �� �h �i �� �i �i �� �i �j �� �j �k �� �k �      �k �� �k 3l �� @l �l �� �l m  � m 1m � �o �o � �o �o � �o �o � �o �o � �o �o � �o �p  � �p �p 0� �p nq 8� pq �q H� �q �q L� �q �q P� �q �q T� �q r X� r �r \� �r �r l� �r t p� t gt |� pt :w �� @w �w �� �w ey �� py �z �� �z �{ �� �{ 7} �� @} �~ �� �~ g�  � p� x� � �� �� � �� ׀ � �� � $� � �� (� �� �� 0�  � ,� <� 0� �� L� �� Q� \� `� � d� �� ,� p� 0� m� t� p� y� �� �� �� �� �� �� �� �� ˆ �� І �� ��  � &� �� 0� :� �� @� ^� �� `� j� �� p� � �� �� �� �� �� �� �� �� �� �� �� ҇ �� �� � �� �� � �� � ň �� Ј �� �� �� T� �� `� � �� �� >� �� @� �� ��  � )�  � 0� � � �� �� � �� ;�  � @� v� ,� �� ː <� А ّ D� �� � \� � �� h� �� Ǖ �� Е r� �� �� �� �� �� �� �� �� [� �� `� � �� �� � ��  � �� ��  � d� �� p� e�  � p� y� � �� �� � �      �� ��  � �� � (� � � 0�  � >� 8� @� K� @� P� Y� D� `� U� H� `� �� T� �� ͞ \� О &� d� 0� �� l� �� � t�  � �� �� �� *� �� 0� �� ��  � �� �� �� �� �� �� ƣ �� У  � ��  � "� �� 0� I� �� P� Z� �� `� �� �� �� �� �� �� �� �� �� ʤ �� Ф ڤ �� � � �� � �� ��  � � �� � �� �� �� � �� � �� � �� ��  � �� � ,� � � 8� � � D�  � )� H� 0� '� L� 0� 5� \� @� ۮ l� � :� x� @� �� �� �� ߯ �� � � ��  � �� �� �� �� �� �� 3� �� @� � ��  � s� �� �� � �� � ų �� г i� �� p� � ��  � �� � �� k� � p� � ,� � � 8�  � �� L� �� �� `� �� ֹ d� � �� h�  � � l�  � � �� � � ��  � �� ȩ �� � �� � �� ��  � �� Щ �� � �� � 0� �� 0� �� �� �� �� T� �� �� �� �� �� |� �� �� x�  � )� ,� 0� ?� (� @� J� �� P� Q� �� `� �� ܫ �� �� ث �� �� 8� �� �� 4� �� �� �      � �� � �� � 4� ܵ @� O� Ե P� U� X� `� a� L� p� �� ̵ �� �� \� �� �� P� �� J� �� P� W� �� `� C� �� P� j� ܪ p� �� ت �� �� Ĭ �� C� �� P� Y� �, `� i� �, p� u� �, �� ,� �, 0� �� @, �� �� ,  � �� h, �� \� , `� }� , �� �� �+ �� � �+ � P� �, P� Y�  . `� i� . p� u� �- �� ,� �- 0� �� t- �� �� D-  � �� �- �� \� L- `� }� <- �� �� �+ �� � �+ � P� �- P� �� �� �� �� �� �� �� 8- �� �� (- �� �� 8+ �� ��  + �� &� �+ 0� D� �+ P� �� H+ �� M� �+ P� �� @+ �� �� 0+ �� �� (+  � ?�  - @� �� �, �� �� �, �� _� �, `� �� + �� �� + �� �� - �� �� l.  � �� \. �� �� <+ �� � `+ � �� h+ �� �� �+ �� M� T+ P� �� �+ �� � �+  � W� �+ `� �� x+ �� �� 4. �� Q� . `� ��  . �� !� . 0� \� + `� w� + �� �� H. �� �� �� �� �� ��  � )� � 0� ?� � @� d� �� p� � �� �� �� x� �� �      �� �� �� �� � �� �� � �� � ��  � O� � P� u� ب �� �� ,� �� �� �� �� �� � �� ��  �� �� (� �� �� �� �� �� � �� ��   � I� P� P� ~� D� �� �� � �� V� 4� `� o� $� p� �� � �� �� � �� !� � 0� A� T� P� �� l� �� �� @� �� �� ȵ �� >� ,� @� H� @� P� X� <� `� �� �� �� �� �� �� �� Ԫ �� �� �� �� �� Ъ �� � � � @� � @� �� � �� �� � �� �� � ��  � ��  � g� �� p� |� �� �� ��  � �� �� �� �� �� � ��  � @�  � N� 8� P� \� <� `� �� L� �� �� (� �� )� � 0� <� $� @� �� 4� �� �� x� �� �� D� �� �� �� �� �� �� �� �� ��  � � T� � � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� L�  � � `� � � @�  � $� �� 0� :� \� @� L� p� P� T� �� `� �� �� �� � ��  � ,� �� 0� a� �� p� x� �� �� �� P� �� �� d� �� �� H� �� ��    � � �� � � ��  � �� h� �� H� P� �      P� H� t� P�   ��    �  T� �  � \� � � X�   + �� 0 B � P X l� ` k h� p t �� � � t� � � $G � � <M � � w � � x� �  ��  � �� � � �� � � �� �   ��   r l� � � |� � � �� � � � � � l� �  ��  j �� p | �� � � �� � � �� � R �� ` l �� p � �� � � �� � � ��    X�   \�   - �� 0 8 �� @ � �� � � � � � 0� � � � � � ,� � 	 <�  	 *	 �� 0	 8	 �� @	 D	 �� P	 T	 � `	 j	 �� p	 |	 �� �	 �	 �� �	 �	 \� �	 ,
 H� 0
 <
 X� @
 p
 h� p
 x
 X� �
 �
 �� �
 �
 �� �
 �
 �� �
 �
 �� �
 �
 P�    `�  r  � � � �� � s 0� � � @�   � � � 5 � @ N �� P { d� � � t� � � �� � � �� � � \� � � �� � � � � 8 ظ @ c ` p � ` � � �_ �  �]   C ` P s �_ � � �      �\ � � �\ � � ` � >  ` @ c �_ p � �] � � �\ � � �\ � � �] �  �]   ) �\ 0 ~ �_ � � �` � � �` � . �` 0 S �] ` � �` � � �` � � �\ � � �\ � . �` 0 ~ �` � � �` � � �] � � �\ � � �\   # �] 0 S �] ` i �\ p � �` � � �� �  ��   n p� p �  � � � �� � � `�    @�   <�   n �� p � x� � � d� �  �   ( 8� 0 9 0� @ c (� p �  � � � 4� � � h�   # l� 0 S h� ` � L� � � � �  d�  3 <� @ H T� P X P� ` � \� � � T�   # @� 0 S 0� ` h L� p y D� � � @� � � 8� � � H� � > D� @ A 8e P d ,e p � 0e � � De �  4e  � Le � M 8� P � @e � � <e � H He P Q �� ` t �� � � �� � � ��      ��    �  ē �  _! p� `! �! �� �! �! �� �! �      X" �� `" Y#   `# Z$ �& `$ q% �m �% �& \m �& �' <� �' �(  � �( �( ,� �( �( �  ) ,) �� 0) \) � `) �) �� �) �* � �* �*  � �* �*  �* |+ �� �+ , �  , �, � �, �- � �- �-  �- �- ��  . . �� . .   . �.  �. �/ �� �/ �/ � �/ �/ L�  0 0 H� 0 0 �  0 �0 �� �0 �0 �  1 n1 �� p1 �1 � �1 N2 �� P2 �2 � �2 �2 �� �2 �2 � �2 N3 �� P3 �3 � �3 .4 �� 04 �4 � �4 5  � 5 ~5 0 �5 �5 (� �5 ^6 8 `6 �6 � �6 >7  @7 K7 0� P7 [7 @ `7 �7 � �7 >8 ( @8 �8 � �8 9    9 ?; � @; �< ��  = �= �� �= �> � �> �@ P  A �B l� �B �C 4� �C �D D �D �E ( �E �F �� �F >G �� @G �G � �G �H T �H �I T� �I .J @� 0J �J � �J �J l� �J �J �/ �J �J 82 �J �J �1 �J �J �1 �J �J 04  K 	K 84 K K �Q  K $K �W 0K 4K $~ @K EK 0� PK UK �0 `K iK �0 pK uK @3 �K �K H3 �K �K <1 �      �K �K D1 �K �K �3 �K �K �3 �K �K � �K �K � �K �K ��  L L �� L L �  L %L � 0L JL �� PL UL Ȅ `L eL ܄ pL uL Ą �L �L ̄ �L �L �� �L �L ؄ �L �L p� �L �L ,� �L QM �� `M �M $�  N qN `� �N �N (� �N $O P� 0O �O � �O �O �� �O �O 0�  P P X� �P �P �  Q ,Q �� 0Q uQ  � �Q ,R \ 0R wR L �R �R �^ �R �S 8' �S �S  � �S (T 0 0T BT 8� PT zU 8� �U �V �� �V ,W H� 0W BW 4� PW �W d� �W PX �� PX �X �� �X �X <� �X %Y l� 0Y �Y �� �Y �Y �� �Y �Y ��  Z Z D�  Z ?[ �� @[ I\ �� P\ |\ � �\ �\ @� �\ ] H�  ] �] � �] �] � �] �] H� �] �^ ��  _ 	` �� ` <` $� @` �` l� �` &a �� 0a Ga H� Pa �a �� �a �a D� �a b $  b 7b � @b �b  �b �b � �b Hc � Pc "d � 0d �d 8 �d �d �^ �d �d �  e e  e .e | 0e 3e   @e �e � �e �e � �e �e | �e 1f p @f Hf l Pf �f � �f �g �      h �g gh � ph �h � �h i � i i �  i �i �  j ;j � @j jj �� pj �m �� �m 	p �� p Ky �� Py �� 8 �� �� �� �� ؃ � �� � , � 3� ( @� ��   �� �� �  � #� $ 0� S� � `� h�  p� x�  �� �  �� _�  `� �� � �� ؆ � �� �  �� ��   � H� � P� �� � �� ��  �� � �  � C�  P� s�  �� � � �� 8� T @� c�  p� �� � �� �� , �� �� ( �� /�  0� �� � �� Ê � Њ � `  � (� $ 0� 9�  @� �� x �� ؋ l �� �   �� _� � `� �� � �� �� � �� /� � 0� x� D �� �� � �� Ӎ � �� � � �� �� �  � o� � p� ߎ � �� � � � X� � `� h� � p� y� � �� ȏ � Џ � �  � )� � 0� �� � �� Ð � А � �  � o� � p� �� 8 �� � � � � �  � (�  0� 8�  @� �� � �� � �  � C� � P� �� h �� ��  �� ��   �� � \ � X� t `� i�  p� �      ߔ � �� �� |�  � � <� � @� T� @� �� @� �� ̕ P� Е  � `�  � � 0� � @� 0� @� �� � �� ̖ ,� Ж ؖ <� �� � Ĉ � � p�  � $� d� 0� `� �� `� �� �� �� ̗ �� З  � ��  � 0� x� 0� �� d� �� �� t� �� � �� � 5� �� @� H� (� P� ]� �� `� h� @� p� ؙ �� �� � �� �  � ��  � � Ȉ � �� ܈  � B� � P� Z� 8� `� e� L� p� t�  � �� �� �� �� �� H� �� �� �� �� �� �� �� � � � ]� �� `� l� � p� �� � �� �� <� �� �� P� �� Μ 0� М G�  � P� T� (� `�  Љ Н !� �� 0� ƞ �� О N� �� P� ͟ �� П �� ĉ �� �� D� �� Ƞ h� Р ߠ x� � �� X�  � � T� � � ��  � <� �� @� K� P� P� �� @� �� ӡ 8� � � <� � !� L� 0� 5� D� @� �� (� �� �  � � c� � p� �� 4� �� ģ ܥ У �� ��  � � x� � @� x� @� �� p� �� �� t� �� Ѥ �� � Y� `� `� �� X� �� � P�  � d� l� p� �� �� �� �� <� �      �� �� ȣ �� ̦ T� Ц ?� ȥ @� D� إ P� �� � �� M� � P� \� � `� �� �� �� �� L� �� Ũ `� Ш Ԩ 4� � � ԥ � �� \�  � 	� �� � � ��  � P� � P� ک  � � � � � !� � 0� 4� P� @� E� d� P� b� D� p� Ȫ ܧ Ъ Ԫ <� � �� �� �� (� �� 0� � ��  � � �� � �� �� �� ï �� Я � X� � � |�  � /� �� 0� F� l� P� [� h� `� h� �� p� �� �� �� Ʊ  б ޱ �� � � � � � � � � �  � B� P P� g� � p� �� �� �� Ƶ   е ޵ �� � � �  � C� �% P� W� �% `� �� 4 �� �� �% �� �� � �� ׸ � � � � � 3� � @� c� � p� �� � �� �� �� �� ù H й ѹ L � � �$ � 	� �$ � <� �$ @� c� �$ p� �� �$ �� �� �$ �� � � � � ,  � � 0 � X� � `� �� � �� �� �  � #� �
 0� S� �
 `� i� 8 p� y� < �� � �
 � _� �
 `� Ͻ �
 н � P  � h� � p� �� � �� � x" � � �      |"  � )�  0� 9�   @� �� �" �� � �"  � �� �" �� �� | �� �� �  � 7� � @� �� �  � _� � `� c� D p� �� � �� 	� � � �� � �� &� h 0� O�  P� K� � P� T� � `� �� � �� ^� � `� t� � �� �� � �� ?� � @� �� � �� �� X# �� [� �' `� �� t' �� � �# � / l# 0 3 ( @ � t# � � �# � ; �# @  D'  [ �# ` �" \' �" �' �# �' �/ �* �/ L2 �' P2 K4 �' P4 �4 d# �4 5 \# 5 o5 |# p5 ZE l `E JU  PU �U t �U +V l 0V X � X \Y � `Y i 8( i �x �' �x +y D  0y �y <  �y k{ �( p{ �| �( �| C} � P} �} � �} ~ �	 ~ .� �	 0� z�  	 ��  � �  � s� `  �� ސ X  �� >� �! @� � �!  � ݛ �  �� �� l  �� �� |�  � �� �� �� � ��  � .� � 0� 3� � @� F� $� P� S�  � `� Ц @� Ц /� � 0� _� � `� n� T� p� v� X� �� �� \� �� �� P� �� �� `� �� � T� � � t�  � �      #� d� 0� �� @�  � N� (� P� � �� � � ��  � Q� �^ `� n� ȯ p� � �^  � C� �g P� W� �g `� ��  ] �� �� �g �� Ӯ ̯ � � h�  � .� ԯ 0� � � � 3� `� @� G� T� P� r� x� �� �� X� �� �� � �� 0� $ 0� D� L P� v� � �� h� � p� ��  �� S dq ` C �p P � �q � C q P �( r �( �1 �r �1 �8 �o  9 _9 d `9 �9 �c �9 : d  : : d �: �: d �: \; �q `; �; �p �; \< r `< �< \q �< \= xr `= �= �r �= �> �r �> �C �p �C �E  p �E �G 0p �G I `p I kI �q pI �I �p �I +J r 0J �J Tq �J �J pr �J KK �r PK #X �) 0X :e �( @e �q �) �q ~ H)  ~ ^� D* `� >� �* @� � � � X� 8� `� (� @� 0� �� ��  � �� �� �� {� � �� � l�  � � �� �� �� t� �� ?� �� @� �� �� �� �� |�  � |� 8� �� �� ��  � |� �� �� �� �  � |� ؠ �� �� 8�  � �� (� �� �� �� �� �� ؞ �� � � � +� �� 0� �� 0� �      �� �� x� �� K� �� P� �� �� �� � Р � k�  � p� �� �k �� � �m � �� n  � L� @n P� =� hn @� �� �k  � S� �n `� �� �n �� � Hd  � [� 0d `� �� 8d �� �� @d �� K� �m P� �� 8n �� � `n � k� �n p� �� @m �� 2� �n @�  �m  X �n ` � �n � � �m   6 0n @ x Xn � � �n �  ��  z x� � ~ �� � �	 � �	 � �   � x� � � D� � � l� � � �� �  ��  N �� P � �� � � ��   [ ܜ ` � � �  <�   \ � ` � ,� � � �� � � d� � A �� P � �� � � Ԝ �  ��  H $� P X �� ` e (� p u � � � xf � � |f � � \f �  Tf   C Xf P g df p � � � � �\ � � �\ � � � � � �� �  Ԕ   C ̔ P s Д � � ܔ � � � � � p� � � t� �  �]  3 �] @ c �] p � 0c � � 4c � � �\ � � �\ � > 8c @ � �      @c � � Hc �   �   3  H� @  c  P� p  �  �� �  �  �� �  �  `� �  �  d� �  >! �� @! �! �� �! �! �� �! " �e " G# |o P# �$ do �$ N& �h P& �& �e �& �& �\ �& ' �e  ' Y* �h `* �, o �, �/ �n �/ �2 4o �2 �G Lo �G %K o 0K �Q �s �Q �S �o �S �U �o �U ?V �e @V �V �e �V �V �e  W #W � 0W �X  � �X KZ � PZ +\ \� 0\ �\ ,� �\ �\ l� �\ �\ 4�  ] �_ D� �_ �b �� �b [e �� `e �h ؝ �h ,| � 0| � �� � �� � �� �� P� �� �� 8� �� � $�  � � � �� ߊ <� �� �� �h �� �� xe  � d� ,k p� A� ,� P� �� � �� �� Й �� �� � �� Ē �A В ג �A �� � xA � �� �A  � � |A � �� �A �� �� tA �� �� �A �� #� �A 0� �� �A �� �� \A �� �� �� �� Ȕ TA Д ؔ XA �� � �B � �� �B  � 	� �B � � �B  � (� �B 0� �� �B �� �� �B �� �� �B �� ו C �� �  C � � �B  � .� �� 0� 8� �B @� H� �B P� �      X� h� `� 2� ,s @� "� �r 0� �� Pb �� � Hb � � �s  � {� ds �� �� x� �� �� @�  � k� Ȑ p� �� �� �� �� � �� ~� �� �� �� lb �� >� db @� ��  m �� �� �l �� �� hl �� d� �k p� �� � �� .� ܐ 0� �� ț �� �� �� �� f� � p� F� �� P� U� 0� `� c�  � p� s� � �� �� (� �� �� 0� �� �� �� �� �� ��  � /� �� 0� �� � �� � �� � �� <  �� *� �� 0� 8� 4� @� g� $� p� ��  � �� �� ,� �� �� (�  � ?� �� @� �� T� �� 3� �� @� H� 4� P� �� $� �� �� � �� �� l� �� �� h� �� �� p�  � � �� � � ��  � (� �� 0� 8� �� @� R� �� `� �� 4� �� � t� � �� �� �� �� � �� � �� � >� �� @� `� �� `� q� 0� �� �� <� �� 	� H� � \� 4� `� �� �� �� �� �� �� �� �� �� (� �� 0� �� �� �� �� ��  � � �  � �� �� �� �� ��  � (� �� 0� � ��  � � H� �� �� �� �� �� �� �� � d� � "� �� 0� p� |� p� �� �� �      �� ��  � �� `� �� `� l� � p� �� �� �� � t� � F� � P� X� � `� �� � �� �� � �� �� ��      ��    G  � P  q  �  �  �  �  �  �  �     �    F �  P q �  � � �  � � �  � � ��   ; �  @ � \  � 
 �   b �  p � �� � 1 �� @ ~ � � � � � � ��   S � ` � `� � � �  �  T    U P� ` � 8� � � ��  	 Y	   `	 �	 $  �	 �	 �  �	 '
 @� 0
 P
 ,� P
 r
 �� �
 �
  �
 �
 4  �
  X�   c �  p � L  � � H� � & @� 0 w �� � �   � 9   @ d �  p � 8� � � $� � � ��   "  0 R ,  ` { <� � � 8� � � �� � � �� � � T�     ��   L l� P y �� � � �� � � �� � � �� � & (� 0 � �E �  `E    �D    ,E  � PE � � �D � ) E 0 y pD � � lD �  E  � �E �  PQ   c @O p � �      �P �  �P  S HP ` � 8N � �  �N  ! C" �N P" �# �M �# �$ �O �$ 3& �O @& �& J �& ) �I  ) �) lJ �) ,+  J 0+ k, �I p, �- <I �- }. �J �. p/  K p/ $0 �G 00 1 (L 1 &2 �L 02 83 �L @3 )4 hL 04 D5 �K P5 K6 xJ P6 �8 � �8 D< h� P< �> H �> �@ �G �@ vA (G �A �D �� �D F �K  F @G DK @G JH dG PH �H �F  I �I 8G �I JJ XG PJ vJ �F �J �J 4G �J �J �F �J K �F  K ;K G @K �K �G  L L G L -L G 0L ML G PL wM �H �M �M �Q �M �M �O �M �M �P �M �M LQ �M �M �P �M #O �H 0O 5O �N @O EO �N PO UO <O `O �P PH �P �P 4N  Q Q �O Q Q DP  Q aR `v pR S �u S �S `t �S �T �t �T �U u �U rV �t �V �W �v �W ?X �u @X �X �u �X Y �u Y pY �u pY �Y Tt �Y �[ �z �[ �] �x �] ` �y ` >b dz @b ^d �w `d ~f Px �f �h (y �h �j �y �j �k �u �k bl t pl �l |u �l ~m Xu �m  n �u  n n t  n �      3n xu @n Xn Tu `n �n �s �n �n �s �n �n <t �n �o �u �o �o @t �o �o Lt �o �o Dt �o �o 0{  p Vq v `q hq $y pq uq \z �q �q �z �q �q `z �q �q Lx �q �q �x �q �q Dx �q �q �x �q r Hx  r (r �x 0r 5r �y @r Er �y Pr or �� pr tr P� �r �r L� �r �r �� �r s ��  s �s �� �s t �� t �t �� �t �t �� �t �t �� �t �t �� �t �t ��  u u ��  u _u H� `u �u � �u Bv \� Pv Xv $� `v �v �� �v �v �� �v �v ,� �v �v (�  w 
w 0� w w l�  w (w T� 0w 8w `� @w Hw d� Pw `w h� `w �w �� �w �w 4�  x {x p� �x �x �� �x �x �� �x y �� y 0y �� 0y Ay �� Py �y �� �y �y � �y ,z �� 0z Pz �� Pz xz �� �z d{ �� p{ �{ d�  | �| x� �| �| �� �| �| �� �| x} �� �} �} � �} �} �� �} �~ l� �~  �  S �� ` o �� p � $� � � �� � � <� � � T�  � P� �� P� �� �� �� ́ �� Ё � ��  � c� 4� p� �� �� �      �� �� �� �� � ��  � ;� |� @� G� T� P� e� �� p� �� �� �� �� �� �� � h�  � � |�  � .� \� 0� S� `� `� s� x� �� �� �� �� Ä �� Є � P� �� +� L� 0� ņ � І � <� �� B� D� P� �� H� �� � @�  � ^� �� `� �� �� �� � x� �� G� �� P� u� � �� Ê �� Њ �� �  � � ��  � f� �� p� �� �� �� � ��  � w� �� �� �� �� �� ό �� Ќ �� � �� � ��  � B� �� P� r� �� �� �� � �� � ��  � &�  � 0� M� �� P� �� � �� � �� �� G� �� P� �� �� �� ֏ �� �� �� ��  �  � �  � B� �� P� r� �� �� �� �� �� ː �� А � �� � � �� � 8� �� @� E� � P� p� x� p� �� ,� �� ȑ �� Б �� ��  � � t� � � ��  � z� �� �� Q� � `� �� � �� �� � �� �� �� �� � �� � X� �_ `� �� �_ �� �� \_  � H� x_ P� �� �_ �� � @_ �  � �  � h� �� p� �� �� И � p`  � g� �` p� �� 8` �� � T` � W� �` `� �� �      ` �� �� �� �� (� �� 0� �� 8� �� � � � 7� D� @� �� ԍ �� ؝ �� �� '� (� 0� |� �� �� �� �� �� �� |�  � b� 0� p� �� � �� �  � � \� �� `� �� ̎ �� �� �  � L� �� P� �� `� �� Ȣ @� Т :� h� @� �� �d �� g� �d p� Ũ pd Ш !� �d 0� �� �d  � U� Td `� z� t^ �� Ԫ `^ � 4� Pe @� �� �� �� �  � � װ p� � 5� � @� �� � �� g� <� p� Ų ̒ в � � � D� ، P� �� ȓ �� � �  � C� �� P� k� �� p� �� �� �� ʴ L� д  � 4�  � >� �� @� a� 8� p� �� � �� ��  � �� � �� � �� ��  � ¶ �� ж � 0�  � S� �� `� �� �� �� b� � p� &� �� 0� 3� �� @� � X� � �� p� �� �� �� �� �� ��  � ǽ �� н � ,� � �� �� �� � t� � [� �� `� =� �� @� f� � p� t� 8� �� �� � �� �� �� �� 8� <� @� �� H� �� �� X� �� 
� t� � � ج �� �� �  � \� d� `� �� �� �� �� Ԭ �� �� D� �� � ��  � �      4� `� @� L� �� P� U� h� `� e� \� p� �� T� �� �� �� �� �� �� �� � t� � [� (� `� r� � �� ��  � �� �� � �� �� P� �� �� �� �� � $� � �� ,� �� �� � �� j� @ p� x� < �� �� �f �� �� 8 �� �� 4 �� �� � �� �� % �� �� d� �� �� l �� &� D 0� Q� �� `� �� �� �� �� ĳ �� �� T� �� �� <� �� � �  � A� з P� m� Գ p� �� d� �� �� D� �� �� � �� � ط � -� ܳ 0� T� l� `� o� H� p� �� d� �� �� `� �� @� �� @� �� p �� `� �� `� �� x �� �� �� �� n� � p� V� � `� +� � 0� w� <� �� �� � �� � l�  � f�  p� �� L� �� � � � W� �� `� �� @ �� �� \�  � O� � P� �� �� �� ��  �� (� � 0� h�   p� �� L� �� �� � �� � � � H� 0 P� �� d� �� �� � �� �� �  � D� P P� �� �� �� �� � �� � $�  � d� X p� �� �� �� �� � �� 6� �� @� �� ( �� �� \� �� � � � V� �� �      `� ��  �� �� T� �� .� � 0� v� �� �� �� 8 �� � |� � N� � P� �� �� �� ��   �� .� �� 0� n� � p� �� �� �� � � � N� t� P� �� � �� �� � �� &� � 0� n� l� p� �� � �� � ,�  � �� h �� �� �� �� P� � P� �� <� �� (� p 0� �� �� �� �� � �� X� D� `� �� x �� 0� �� 0� �� � �� �� 4�  � h� ` p� �� �� �� 0� � 0� d� D� p� �� � �� �� <� �� �� � �� � X� � �   � <� �� @� N� 4 P� �� � �� ^� � `� �� 4� �� n� � p� �� �� �� �� ` �� �� �� �� �� d �� �� p� �� �� ( �� � t� � /� , 0� �� x� �� d� 0 p� 
� �� � �� T �� �� �� �� �� h �� �� �� �� �� l �� �� �� �� $ � 0 X $� `  �  Z � ` <	 � @	 � �� � l x p S �� ` � h � � P� � �  � * � 0 b � p z t� � � d� � � T0   r �/ � � @/ �  D/   �/   � �      �/ � � �/   3 �/ @ 9 06 @ H @6 P [  �/ `  �  �. �  �! D4 �! �# H0 �# $ p. $ C&  / P& ~'  / �' 4( 0 @( * $0 * �* 80 �* �, 0 �, �- �. �- . �. �. �3 �. �3 E5 �/ P5 �6 l/ �6 58 �/ @8 �9 H/ �9 �9 D9 �9 : �4  : \: �4 `: �; �5 �; K< �2 P< �< `2 �< = �1 = W= �1 `= a> l2 p> �? H2 �? K@ @2 P@ e@ <2 p@ �@ �. �@ �A < �A �A  < �A �C (2 �C �C �. �C �D $: �D 
G �2 G mG |. pG sI 0/ �I �J / �J tK �2 �K MM �2 PM �M �2  N �O �2  P AQ �. PQ �Q �.  R W �.  W �X 2 �X Z �1  Z �[ 2 �[ ] �1  ] d] $? p] �] p: �] �] `: �] o_ �; p_ �_ l6 �_ ` T6 ` �` �1 �` 
a �8 a a �1  a �b p1 �b d t6  d �e �6 �e �f �5 �f ]h H1 `h �i �6 �i k  7  k 8l T5 @l �l �9 �l �m 49 �m =n �9 @n o �5 o Wo L< `o �o 4< �o rp 4 �p �p �> �p �p 44 �p >r �3 @r �s T< �s Vu �< `u �      �v h; �v x �3 x my �< py �z  = �z �{ 4; �{ �| �? �| 9} ? @} �} t? �} �~ �; �~ � `\ � T� PZ `� �� �[ �� � \  � D� X[ P� �� HY �� � �Y �� 4� �Y @� �� �X �� ԋ �Z �� $�  [ 0� ~� �T �� ُ �T �� &� 4U 0� � �T � %� <T 0� Q� �S `� N� �U P� @� �U @� �� `R  � ܗ �V �� �� dW  � � �W � ��  W  � #� �V 0� 0� @U 0� �� 8� �� 
� �� � � �R � � xR � ^� �Q `� �� ,� �� � TV � !� V 0� B� $R P� � �Q � �� �Q �� [� R `� �� �Q �� �� �Q �� �� �F  � )� �F 0� K� �Q P� 	� HR � � �Q  � =� �Q @� ]� �Q `� �� �S �� �� �\ �� �� �Z �� �� \ �� ų \\ г ճ �[ � 3� dS @� E� �Y P� U� �Y `� e� LZ p�  � S  � � DY � � �Z  � %� T[ 0� �� |} �� )� �| 0� � |{ � ݺ �{ � �� 4| �� �� �{ �� � �} � _� �| `� Ͼ �| о 0� } 0� �� } �� ۿ p{ � �� � �� � � �� O� @� �      P� /� �� 0� �� <  � �� � �� �� x� �� o� ܀ p� m� �| p� � 8{  � �� �| �� 5� t| @� �� �| �� �� 4{ �� � �| � (� p| 0� f� �s p� �� �s �� �� X{ �� d� �| p� s� \{ �� �� h{ �� �� `{ �� �� t� �� &� ,} 0� 8� t� @� E� �� P� i� � p� y� �� �� �� � �� �� � �� �� � �� �� � �� �� � �� �� �  � � ؀ � � <�  � �� �� �� o� �� p� �� � �� � �� � +� Ĵ 0� h� � p� �� |� �� �� t� �� �� д  � G� \6 P� �� D6 �� `� �0 `� �� �8 �� �� �0 �� � �0 � ^� �7 `� �� �8 �� �� �4 �� �� X0 �� �� �7 �� �� @8 �� D� �4 P� �� �9 �� g� $9 p� �� �8 �� �� �5 �� � << � Z� $< `� "� (3 0� j� �> p� y� D3 �� �� �2 �� 2� �= @� �� �> �� �� �: �� �� �2 �� �� `= �� ��  > �� D� �: P� �� �? �� g� ? p� �� �> �� �� �; �� v� �F �� �� dF �� �� �E �� �� 0F �� �� TF �� 0� �E 0� �� F �� � �      |D  � U� xD `� �� F �� i� �F p� �� d6 �� 
� L6 � �� $1 �� �� �8  � 	� @1 � K� �0 P� �� �7 �� �� l8 �� �  $5 �  � �0 � � T7 � � 8 � / �4 0 � �9 � ? 9 @ �  9 � d 6 p � D< � 
 ,<  � �3 � 
 �>   �3   c	 t3 p	 �
 �= �
  L>   ;  � L3   � 4= � � �= � o �: p � �?    �> � � �> � � �; � H g P � h � � hg � ( �f 0 � @ � h @g p � �^ � � |^ � � �g � X �� ` � D%   � �� � 8 h� @ � % � x �� � � �� � � � � � � � � $h � � th � h �g p H Lh P � P^ � � @^ � � �h � � �� � �  � �  x! t� �! X" Ė `" �" Ȍ �" �" �� �" �" � �" # @�  # A# � P# m# � p# �# �� �# �# �� �# �# ��  $ Q$ �� `$ e$  � p$ u$ $� �$ �$  � �$ �$ � �$ F% 8� P% S% Ȃ `% h% �� p% q% �� �% �      �% � �% �% Ѓ �% �% ԃ �% & ��  & '& � 0& |& H� �& �& ȃ �& �& ��  ' �' �� �' +( � 0( ) P� ) �) � �) �) �� �) �) ��  * * Ă  * ]* ܃ `* �* �� �* �* ؂ �* + |� + + Ԃ  + C+ �� P+ S+ ̂ `+ �+ ؃ �+ �+ Ђ �+ �+ ,�  , C, � P, �, (� �, �, � �, - �  - 3-  � @- S- x� `- �- 0� �- �- |�  . Q. �� `. h. � p. x. �� �. �. Ԅ �. �. � �. F/ � P/ S/ � `/ k/ Є p/ q/ ܂ �/ �/ � �/ �/ �� �/ �/ �� �/ 0 �� 0 0 ��  0 m0 @� p0 �0 �� �0 �0 ��  1 �1 �� �1 2 �  2 �2 d�  3 �3 ,� �3 �3 �� �3 �3 � �3 4 � 4 P4 �� P4 |4 �� �4 �4 �� �4 �4 P�  5 5 �� 5 35 x� @5 C5 �� P5 �5 �� �5 �5 � �5 �5  � �5 36 �� @6 �6 �� �6 �6 �� �6 7 � 7 #7 � 07 C7 L� P7 �7 � �7 J8 �f P8 X8 �f `8 
9 �f 9 9 �f  9 P9 0^ P9 x9  ^ �9 �9 �f �9 Z: $� `: h: P� p: ; ��  ; (; L� �      0; `; �� `; �; �� �; �; T� �; �< xc �< y= �c �= Y> Pc `> 9? �c @? d? H] p? ? �\ �? �? �c �? i@ � p@ IA @� PA )B ȑ 0B 	C � C 4C �� @C OC h� PC _C h� `C vC �e �C �C �e �C �C �e �C �C �e �C D �] D D $]  D /D �e 0D FD L� PD fD T� pD �D H� �D �D P� �D �D �� �D �D �� �D �D X�  E E �e  E :E p @E VE �e `E vE �e �E �E l �E �E �e �E �E x] �E �E  ]  F F �e F &F  � 0F JF L# PF fF � pF �F �� �F �F H# �F �F � �F �F ��  G G �� G G �  G AG H� PG qG � �G �G � �G �G �� �G �G �� �G �K i �K 'L |b 0L �L xb �L �L H� �L M @�  M rM �b �M hQ �� pQ �Q �� �Q (R � 0R `R l� `R �R d� �R S ��  S AS � PS qS ȷ �S �S ̳ �S �S \� �S �S @� �S �U he �U �W de �W X `] X X ]  X /X le 0X (Z �� 0Z (\ ܓ 0\ T\ ؋ `\ o\ �� p\ \ � �\ \]  a `] <^ pa @^ _ �`  _ �_ �      Ha  ` $` (] 0` ?` �\ @` O` �a P` ,a �a 0a b b b �b �a �b �c �a �c �c 0]  d d �\ d d <b  d �d ��  e �e � �e �f p� �f �g �� �g �g �� �g �g X� �g �g � �g �h <� �h �i �� �i �j � �j lk d� pk �k �� �k �k \� �k �k �� �k �p hj �p q $_  q �q  _ �q �q @� �q -r 8� 0r �r (_ �r mw �i pw �w 4_ �w cx 0_ px �x � �x �x �  y ]y 8_ `y �~ �� �~ 4 �� @ � �� � � �� � M� �� P� �� �� �� � 0� � �� �� �� � �� � @� d� @� �� \� �� �� ��  � $� �� 0� ?� `� @� d� t� p� � P� �� �� �� �� �� �� �� � �� �� �� ��  � $� �� 0� ?� d� @� d� |� p� � T� �� �� �� �� �� �� �� � �� �� �� ��  � $� �� 0� ?� h� @� d� �� p� � X� �� �� �� �� �� �� �� Ŋ ̸ Њ ъ ȸ �� � и �� �� Ը  � �� (m �� �� Л �� ��   �� >�  @� ��  �� ڐ T �� � $  � �� � �� � � � k� � p� �      �� \ �� � 4 � K� �� P� �� |� �� ѓ L� �� ͙ �� Й �� � �� �� |� �� Σ �� У � h�  � _� p� `� �� ��  � �� �� �� �� `� з ط \� � � T� � � H�  � [� 8� `� v� �� �� �� D� �� �� L� �� �� �� �� �� �� �� �� �� й �� ��  � � �� � � ��  � պ �� � 	� �� � d� �� p� ż � м � �  � g� � p� �� ` �� � | � W� � `� �� D �� � p� � (� P� 0� �� � �� �� � �� '� � 0� |� L �� �� h �� � �  � l� 0 p� �� 4� �� �� � �� V� �� `� �� h �� �� �  � L� 0 P� �� L �� �� � �� <�  @� p� �� p� �� �� �� &� �� 0� x� T �� �� � �� �   � h� 8 p� �� p �� �   � @� �� @� �� �� �� �� L� �� �� H� �� ^� t� `� � �� �� �� 4� �� �� � �� ��  � �� �� � �� �� �� �� [� P� `� �� d�  � �� P� �� _� �� `� � x�  � %� ,� 0� <� 8� @� [� �� `� {� �� �� �� �� �      �� �� �� �� 	� l� � /� � 0� 4� `� @� I� \� P� u� �� �� �� $� �� �� �� �� �� 4� �� �� �� �� �� � �� �� �� �� �� ��  � T� � `� �� � �� �� (� �� O� �� P� T� �� `� �� �� �� �� �� �� �� p� �� 3� x� @� w� �� �� �� $� �� J� �� P� �� �� �� �� �� �� �� ؆ �� � ��  � @� �� @� `� 8� `� �� P� �� �� h� �� $� 0� 0� f� D� p� �� 4� �� �� H�  � <� ԇ @� �� ̇ �� �� �  � @� H� @� �� <� �� �� ,� �� �� 4� �� �� ,� �� ��  �  � � ��  � ;� �� @� ��  � �� �� �  � V� � `� �� T� �� 6� �� @� �� � �� �� (� �� I� � P� i� d� p� �� �� �� A� `� P� �� |� �� �� X�  � V� P� `� �� t� �� � ��  � 9� p� @� �� 8� �� �� �� �� :� ܇ @� �� � �� � \�  � +� \� 0� �� ȅ �� �� � �� :� d� @� �� �� �� ]� @� `� e� $� p� �� �� �� �� �� �� I� Ȇ P� �� �� ��  � ��  � ?� � @� R� � `� t� �      �� �� �� �� �� �� t� �� � Ȋ � \� ؊ `� �� � �� �� � �� �� ؅ ��  � �  � � `� � � �  � /� �� 0� {� � �� �� � �� � ��  � 2� �� @� T� ܅ `� |� �� �� �� p� �� �� �� �� <� Њ @� �� �� �� �� � �� �� ԅ �� �� � �� �� \� �� �� �  � � �� � %�  � 0� E� �� P� �� � �� !� �� 0� F� � P� x� �� �� �� @� �� �� �� �� � �� � � t�  � W� �� `� �� �� �� �� `� �� � \� � �� �� �� �� ��  � � H� � � ̦  � $� Ħ 0� 4� Ȧ @� D� �� P� �� d� �� Q� (� `� �� � �� �� x� �� A� <� P� U� @� `� n� L� p� �� �� �� �� �� �� �� ��  � '� �� 0� y� �� �� �� (� �� �� t� �� �� p� �� �� ��  � � 8� � � ģ  � *� H� 0� 1� Х @� D� 0� P� a� �� p� �� � �� �� �  � -� �� 0� �� �� �� �� �  � � �� � X� �� `� �� �� �� �� �� �� �� �� �� ' 	 �� 0 	 Q 	 <� ` 	 � 	 �� � 	 !	 Ĥ 0	 �      L	 �� P	 f	 � p	 �	 �� �	 �	 �� �	  	 P�  	 9	 h� @	 v	 �� �	 �	 8� �	 		 �� 	 4	 �� @	 �	 P� �	 �	 � �	  	 �  	 �	 � �	 �	 `� �	 )	 �� 0	 B	 @� P	 X	 L� `	 �	 D� �	 �	 4� �	 �	 �� �	 	 ��  	 �	 @� �	 �	  �  	 \	 �� `	 �	 l� �	 B	 (� P	 �	 � �	 		 H� 		 o		 0� p		 �		 |� �		 �		 �  
	 w
	 ز �
	 �
	 �� �
	 ?	 в @	 �	 Ȳ �	 	 � 	 r	 �� �	 �	 � �	 	 \� 	 M	 Ф P	 �	 �� �	 &	 � 0	 x	 t� �	 �	 p� �	 �	 ܢ  	 	 $�  	 �	 |� �	 h	 �� p	 �	 T� �	 �	 8� �	 ,	 Ģ 0	 U	 �� `	 �	 ܣ �	 	 �  	 �	 � �	 �	 ħ �	 �	 ��  	 	 ��  	 =	 L� @	 ]	 8� `	 �	 �� �	 �	 ��  	 L	 �� P	 m	 Ч p	 �	 � �	 �	 �� �	 �	 $� �	 �	 ا �	 �	 t� �	 	  �  	 �	 � �	 �	 �� �	 �	 ��  	 	 �  	 =	 H� @	 ]	 4� `	 �	 �� �	 �	 ��  	 L	 �� P	 m	 ̧ p	 �	 � �	 �	 �� �	 �	  � �	 �	 ԧ �      �	 �	 p� �	 �	 � �	 	 � 	 �	  � �	 �	 ؤ �	 �	 �  	 (	 �� 0	 Y	 X� `	 h	 �� p	 �	 �� �	 �	 �� �	 	 �� 	 {	 ̣ �	 X	   `	 8	 p @	 	 �  	 �	 H   	 0 	  0 	 X 	 � ` 	 � 	 � � 	 h!	 �% p!	 H"	 L& P"	 (#	 �% 0#	 $	 $& $	 @$	 � @$	 h$	 � p$	 �$	 t& �$	 J%	 � P%	 X%	 ( `%	 
&	 � &	 &	 $  &	 P&	 � P&	 x&	 � �&	 �&	 , �&	 Z'	 �$ `'	 h'	 % p'	 (	 �$  (	 ((	  % 0(	 `(	 � `(	 �(	 � �(	 �(	 % �(	 �)	 �
 �)	 y*	 @ �*	 Y+	 �
 `+	 9,	  @,	 d,	 � p,	 ,	 @ �,	 �,	 h �,	 i-	 �" p-	 I.	 # P.	 )/	 �" 0/	 	0	 �" 0	 40	 h @0	 O0	 $ P0	 _0	 D# `0	 v0	 ( �0	 �0	 0 �0	 �0	 $ �0	 �0	 , �0	 1	 � 1	 1	 `  1	 /1	 4 01	 F1	 $ P1	 f1	 $ p1	 �1	  $ �1	 �1	 $ �1	 �1	 x �1	 �1	 D �1	 �1	 $  2	 �2	 D �2	 �3	 � �3	 �4	  �4	 |5	 l �5	 �5	 d �5	 �5	 0 �5	 �5	 � �5	 �6	 � �6	 �7	 8 �7	 l8	 � p8	 L9	  P9	 t9	 l �9	 �9	 4 �9	 �9	 ` �9	 |:	  �:	 \;	 �      d `;	 <<	 � @<	 =	 <  =	 D=	 H P=	 _=	  `=	 o=	 � p=	 L>	 � P>	 ,?	   0?	 @	 � @	 �@	 � �@	 A	 P  A	 /A	  0A	 ?A	 0  @A	 vA	 � �A	 �A	 � �A	 B	 � B	 RB	 � `B	 �B	 � �B	 �B	 � �B	 �B	 � �B	 &C	 �% 0C	 rC	 �% �C	 �C	 �% �C	 D	 l% D	 @D	 � @D	 hD	 � pD	 �D	 �% �D	 �D	 � �D	 2E	 T @E	 �E	 p �E	 �E	 8 �E	 F	 � F	 8F	 � @F	 hF	 � pF	 �F	 h$ �F	 G	 0$ G	 RG	 L$ `G	 �G	 $ �G	 �G	 � �G	 H	 � H	 8H	 �$ @H	 oI	 �� pI	 �I	 H
 �I	 J	 �
 J	 YJ	 
 `J	 �J	 ,
 �J	 �J	 d
  K	 IK	 �	 PK	 �K	 �� �K	 �K	 �� �K	 �L	 �� �L	 %M	 $" 0M	 wM	 \" �M	 �M	 �! �M	 N	 "  N	 gN	 @" pN	 �N	 �! �N	 �N	 $� �N	 8O	 � @O	 VO	 x `O	 vO	 t �O	 �O	 � �O	 �O	 \ �O	 �O	 � �O	 �O	 T# �O	 P	 P# P	 4P	 p @P	 OP	 @ PP	 _P	 �# `P	 vP	 h �P	 �P	 d �P	 �P	 t �P	 �P	 T �P	 �P	 | �P	 Q	 8  Q	 &Q	 4  0Q	 TQ	 X `Q	 oQ	 8 pQ	 Q	 L  �Q	 �Q	 � �Q	 �Q	 � �Q	 �Q	 | �Q	 �Q	 X  R	 R	 � R	 &R	 T  0R	 �      FR	 P  PR	 tR	 ` �R	 �R	 < �R	 �R	 h  �R	 �R	 �� �R	 �R	 \� �R	 S	 l� S	 S	 L�  S	 VS	 �� `S	 �S	 � �S	 �S	 �� �S	 :T	 h� @T	 vT	  � �T	 �T	 � �T	  U	 Į  U	 ZU	 �� `U	 �U	 �g �U	 �U	 �g �U	 &V	 �g 0V	 rV	 �g �V	 �V	 ^ �V	 �V	  ^ �V	 W	 �g W	 FW	 L� PW	 �W	 (� �W	 �W	 D� �W	 "X	 � 0X	 `X	 �� `X	 �X	 x� �X	 �X	 d� �X	 �X	 �c �X	 �X	 �c  Y	 $Y	 P] 0Y	 ?Y	 ] @Y	 OY	 $d PY	 fY	 p� pY	 �Y	 l� �Y	 �Y	 ȋ �Y	 �Y	 �� �Y	 �Y	 �� �Y	 �Y	 ,d  Z	 Z	 (d  Z	 DZ	 X] PZ	 _Z	 ] `Z	 oZ	 Pd pZ	 �Z	 �� �Z	 �Z	 �� �Z	 �Z	 Ћ �Z	 �Z	 �� �Z	 �Z	 Ȓ  [	 )[	 � 0[	 ?[	  � @[	 �\	 �C �\	 7_	 l� @_	 �_	 D �_	 �_	 �C �_	 !`	 4D 0`	 �g	 �� �g	 ph	 L� ph	 �h	 � �h	 �h	 �C �h	 ,i	 د 0i	 `j	 PD `j	  l	 `D  l	 on	 �� pn	 q	 T� q	 �s	 �� �s	 t	 � t	 t	 �  t	 ht	 <� pt	 �t	 4� �t	 �t	 ,� �t	 au	 �C pu	 �u	 HD �u	 �u	 @D �u	 2v	 8f @v	 �v	  f �v	 �v	 f �v	 "w	 �e 0w	 `w	 �] `w	 �w	 �] �w	 �w	 hf �w	 x	 �� x	 Rx	 x� `x	 �x	 �� �      �x	 �x	 \�  y	 0y	 h� 0y	 Xy	 X� `y	 �y	 �� �y	 �z	 �� �z	 {	 �b {	 W{	 c `{	 �{	 �b �{	 �{	 �b  |	 G|	 �b P|	 �|	 �b �|	 �|	 �� �|	 }	 ��  }	 +~	 �� 0~	 u~	 T� �~	 �~	 �� �~	 	 �  	 e	 8� p	 �	 p� �	 	�	  � �	 @�	 �� @�	 ��	 �� ��	 ��	 �e ��	 ƀ	 �e Ѐ	 �	 p]  �	 �	 ] �	 �	 �e  �	 6�	 � @�	 V�	 � `�	 ��	 � ��	 ��	 �� ��	 ��	 D� ��	 Ɓ	 te Ё	 �	 pe ��	 �	 h]  �	 /�	 ] 0�	 ?�	 �e @�	 V�	 � `�	 v�	 � ��	 ��	 �� ��	 ��	 �� ��	 ς	 �� Ђ	 ��	 ��  �	 �	 � �	 �	 �A  �	 7�	 lA @�	 ̓	 �A Ѓ	 ߃	 �A ��	 s�	 �A ��	 Ԅ	 ,B ��	 E�	 �B P�	 ��	 pB ��	 F�	 |B P�	 ��	 `A ��	 >�	 B @�	 u�	 �A ��	 �	 �A �	 �	 hA  �	 (�	 �A 0�	 ��	 TB ��	 �	 �A  �	 ��	 8B ��	 �	 �A �	 4�	 DA @�	 O�	 <A P�	 _�	 �A `�	 k�	 �B p�	 ��	 �B ��	 �	 $C  �	 /�	 �B 0�	 ��	 �B ��	 ��	 hC  �	 f�	 �C p�	 ֎	 �C ��	 h�	 �C p�	 ��	 �B ��	 ^�	 @C `�	 ��	 �B ��	 Ē	 0C В	 ؒ	 �B ��	 �	  C �	 y�	 �C ��	 �	 C �	 y�	 tC ��	 �	 �      C �	 �	 LA  �	 /�	 @A 0�	 ?�	 �B @�	 J�	 p� P�	 Q�	 `� `�	 v�	 Db ��	 ��	 @b ��	 ĕ	 8] Е	 ߕ	 ] ��	 �	 Xb �	 �	 �� �	 &�	 �� 0�	 T�	 �� `�	 o�	 |� p�	 �	 А ��	 ��	 `b ��	 ��	 \b ��	 �	 @] �	 ��	 ]  �	 �	 tb �	 &�	 ؐ 0�	 F�	 Ԑ P�	 t�	 �� ��	 ��	 �� ��	 ��	 � ��	 ��	 $� ��	 ��	 � ��	 ԗ	 �� ��	 ��	 Lm ��	 ^�	 Tm `�	 �	 �  �	 �	 ��  �	 �	 �� �	 �	 ��  �	 ��	 �k ��	 0�	 h� 0�	 =�	 ح @�	 \�	 � `�	 g�	 �� p�	 {�	 �� ��	 ��	 �� ��	 ��	 �� ��	 ��	 �� ��	 ��	 $ ��	 ~�	 @w ��	 5�	 X~ @�	 s�	 @ ��	 ��	 D� ��	 ��	 � ��	 �	 @  �	 *�	 � 0�	 <�	 �� @�	 N�	 L� P�	 ��	 @ ��	 ��	 P� ��	 �	 <�  �	 k�	 @ p�	 ��	 �@ ��	 Ѯ	 X� �	 +�	 8@ 0�	 {�	 p@ ��	 ˯	 �@ Я	 t�	 �� ��	 ��	 � ��	 ��	 (� ��	 Ʋ	 p� в	 �	 �? �	 [�	 �@ `�	 ��	 A ��	 J�	 � P�	 ��	 d� ��	 ��	  A  �	 �	 t� �	 [�	 T@ `�	 �	 �@  �	 �	 @M �	 �	 �W �	 `�	 w `�	 ��	 (~ ��	 ��	 w ��	 Ǹ	 0~ и	 ո	 w �	 �	 4~ �	 �	 �D  �	 �      �	 �E �	 a�	 � p�	 ��	 �& й	 !�	 � 0�	 ��	 �& ��	 �	  �	 A�	 �& P�	 ��	 � ��	 �	 �& �	 a�	  p�	 ��	 �& м	 !�	  0�	 ��	 �& ��	 �	   �	 A�	 �& P�	 ��	 �k ��	 �	 0� �	 a�	 �k p�	 ��	 H� п	 !�	 \k 0�	 ��	  � ��	 ��	 dk ��	 A�	 � P�	 ��	 lk ��	 �	 � �	 a�	 �k p�	 ��	 (� ��	 !�	 |k 0�	 ��	  � ��	 ��	 �k ��	 A�	 `� P�	 ��	 tk ��	 �	 � �	 a�	 �k p�	 ��	 X� ��	 !�	 �k 0�	 ��	 P� ��	 ��	 �k ��	 A�	 @� P�	 ��	 �k ��	 �	 8� �	 $�	 �� 0�	 ��	 � ��	 ��	 � ��	 F�	 �& P�	 ��	 �& ��	 �	 � �	 f�	 �& p�	 ��	 � ��	 &�	 �& 0�	 ��	 � ��	 ��	 �& ��	 F�	 � P�	 ��	 �& ��	 �	 � �	 f�	 �& p�	 ��	 � ��	 &�	 �& 0�	 ��	 `j ��	 ��	 �i ��	 F�	 � P�	 ��	 (� ��	 �	 $k �	 f�	 ș p�	 ��	 �h ��	 &�	 $� 0�	 ��	 �h ��	 ��	 t� ��	 F�	 i P�	 ��	 |� ��	 �	 �i �	 f�	  � p�	 ��	 �i ��	 &�	 � 0�	 ��	 Tk ��	 ��	 �� ��	 F�	 i P�	 ��	 �� ��	 �	 Lk �	 f�	 � p�	 ��	 Dk ��	 &�	 � 0�	 ��	 k ��	 ��	 �� ��	 F�	 k �      P�	 ��	 �� ��	  �	 �w  �	 P�	 �w P�	 ��	 �w ��	 ��	 �w ��	 ��	 �w ��	 ��	 �w  �	 �	 ,w  �	 3�	 8w @�	 T�	 0w `�	 s�	 <w ��	 ��	 4w ��	 >�	 w @�	 ��	 �~ ��	 �	 �~  �	 >�	 �~ @�	 R�	 D~ `�	 s�	 P~ ��	 ��	 H~ ��	 ��	 T~ ��	 ��	 L~  �	 W�	 8~ `�	 ��	 �~ ��	 S�	 � `�	 ��	 �� ��	 A�	 0� P�	 ��	 � ��	 L�	 h� P�	 ��	 D� ��	 u�	 Ц ��	 ��	 P� ��	 b�	 �� p�	 �	 X� �	 |�	 �� ��	 �	 ��  �	 %�	 �M 0�	 5�	 �M @�	 E�	 �M P�	 U�	 �M `�	 ��	 �� ��	 ��	 `M ��	 ��	 �M ��	 ��	 �M ��	 ��	 �M ��	 �	 �M �	 J�	 �M P�	 ��	 �M ��	 W�	 dX `�	 a�	 X p�	 ��	 �X ��	 ��	 �X ��	 ��	 �X ��	 ��	 �X ��	 *�	 �X 0�	 ��	 �X ��	 ��	 �D ��	 �	 �D  �	 ��	 �9 ��	 j�	 �9 p�	 �	 �?  �	 ��	 T? ��	 
�	 �D �	 D�	 �D P�	 ��	 �D ��	 ��	 �D ��	 6�	 �F @�	 p�	 �F p�	 ��	 t ��	 ��	  t ��	 ��	 : ��	 1�	 t9 @�	 ��	 �? ��	 ��	 4? ��	 ��	 �F ��	  �	 �F  �	 ^�	 t `�	 ��	 t ��	 &�	 �9 0�	 ��	 d9 ��	 V�	 �? `�	 ��	 d? ��	 A�	 �D P�	 ��	 �D ��	 �	 �9  �	 ��	 �      T9 ��	 >�	 �? @�	 ��	 D? ��	 .�	 <4 0�	 ��	 : ��	 ��	 h� ��	 ��	 `� ��	 ��	 d� ��	 ��	 �� ��	 ��	 ī ��	 M�	 �� P�	 ��	 � ��	 ��	  �   
 V 
 � ` 
 � 
 $� � 
 � 
 ,� � 
 ]
 @� `
 �
 �� �
 �
 � �
 �
 �� �
 �
 Ы  
 ~
 H� �
 �
 � �
 �
 �� �
 �
 <� �
 �
 ��  
 
 �� 
 �
 @� �
 0
 � 0
 �
 x�  
 X
 �� `
 �
 ȫ �
 �
 Ȫ �
 S
 �� `
 �
 4� �
 �	
 l� �	
 �	
 L� �	
 �	
 �� �	
 �	
 �� �	
 �	
 |�  

 

 ص  

 !

 T� 0

 1

 �� @

 �

 | �

 Q
 + `
 !
 �s 0
 �
 0�  
 q
 � �
 �
 �� �
 �
 � �
 �
 ػ �
 	
  � 
 
 p�                                                                                                                                                                                                                                                                                                                                                 B   b    0`pP��	 B  �     �      �  �  �  �  	 B  �     �  �  �  �   B        2P  2P  2P  2P  2P  2P  2P   2
0	`pP���	
 ��cG�  �� �� �� �� ��  �	� �
� �� �� �  �  �  �  �  �  �  �    B  �	
 ��'An{         R0`p�	
 ��,  ��� �  �                           20    20 B  �	
 ��8?H              	 b0`
p	P����  �	
 ����� �   �0`pP  �	
 ��U�e��    }     B   B      B0`  �	
 ��)A��������                20 20
 
20`pP��	
 ��S���� �          	 B0`
p	P����  �	
 ��aTf  ���  �����  �������� �������  �                B   20`p R0`p�	
 ��%!+  �� ���� ���@          �	
 ��  20�	
 ��9c u   B  	 �0`
p	P����  �	
 ��un�B��� �i��� ���� ����      ������ �i��� ���� ���������    }      B   20 20`p�	
 ��.�SG����        B   �0`pP  �	
 ��%  O� ��  ���           20 20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 B0`  �	
 ��	 *   20 B0`  �	
 ��	 *   20 B0`  �	
 ��	 *   20 B0`  �	
 ��	 *      20 20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 B0`  �	
 ��#4 /  B   �      B0`  �	
 ��	 *   20 B0`  �	
 ��	 *   20 B0`  �	
 ��	 *   20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   20 B0`  �	
 ��#4 /  B   B0`  �	
 ��	 *   0`                                                                20 20 20 20 20 20 20 20          20    20    20       b0`      20`p b   �   �   �   �   b0`   20
 
r0`pP�
 
r0`pP� 20`p r0 r0 B0`pP   R0 R0 0   r0 R0`p R0`p   
 
R0`pP�
 
R0`pP� R0`p R0 R0
 
R0`pP� R0 R0 R0 R0 B0`pP��   �   �   �   �   b0`pP   20`p �   �   r0 R0`p R0	 B0`
p	P����  �	
 ��:M�
 �� �� �� �  �� ��
 ��
 ��
 �	�    	 b0`
p	P����  �	
 �      ��\)  T�	 |T  ��	 �  ��	 ��  ��	 �  ��	 �T  ��	 �  ��	 ��  ��	 �	   r
0	`pP���	
 ��   ��� �   b   �0 �0 �0 �0 �0   	 	 0` �0    b   b   �0 �0 �0 �0 �0     0   �0    b  
 x
  0`pP�а	
 ��
Ki� �    
 x
  0`pP�а	
 ��
Kj� �     �0`  �	
 ��($q lq �      �0`  �	
 ��($q lq �     	 	 0`�	
 ��O$� �� �  	 	 0`�	
 ��O$� �� �   b   b   20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20�	
 ��  20 20 20 20�	
 ��  20 20 20 20 20 20 20 20 20 20�	
 ��  20�	
 ��  h  0`pP�	
 ���� �� �� �� �       0`pP�а	
 ���� �� �� �� �        
 
R0`pP��	
 ��$B  e� �  �� �         �� �   b0`pP��  �	
 ��0D  i� �  �� �  �� �#  �� ��        b0`  �	
 ��  +{ �      b0`  �	
 ��  +{ �     
 
R0`pP��	
 ��0S  v� �  �� �  �� �  �� ��  
 
R0`pP��	
 ��0S  v� �  �� �  �� �  �� ��   b0`pP��  �	
 ��BU  z� �  �� �  �� �  �� ��  �� �� ��    b0`pP��  �	
 ��BU  z� �  �� �  �� �  �� ��  �� �� ��    r0`p�	
 ��   6p �      r0`p�	
 ��   6p �     
 
�0`pP��	
 ��5  ^� m� �   
 
�0`pP��	
 ��5  ^� m� �                �0 �0 x  0`
p	P����	
 ���:  �� �   x
 h	  0`pP�а	
 ���D  ��� �     
 x  0`pP�а	
 ��o  �� �A   
 x  0`pP�а	
 ��o  �� �A    20`p�	
 ����  �� �h  �� �� �?  �� �  �� ��  �� �� ��  �	� �	� �
  �
�       �
i  �� �� ��  �� �� ��  �� �� ��                     B   B                                                                                    B         20    B   B            2
0	`pP���    20`p B0`   B0`pP      20`p   
 
20`pP�    20`p    B0`pP      20`p   
 
20`pP�    20`p    B0`pP      20`p    B0`   B0`   B0`   B0`pP  
 
20`pP� B0`                              20	 b0`
p	P����   20    B0`   20 B0`   20 B0`   20 B0`   B0`      20 B0`   B0`   B0`pP   b   R0 b   b0`   B      b   B0`pP   b0`   20 B   B0`   B0`      b0`pP      B   20`p    B   20`p R0 R0 20 20       20 20 R0 R0             B0`   r0 B  �	
 ��"-       B0`pP      B0`pP   20`p    B0`   B0`      B0`pP   20 B      B0`pP   B0`pP      R0 R0 b0`     
 
R0`pP��	
 ��*  ?k �      b0`pP  �	
 ��  2!_ t   b0`  �	
 ��-O H$   20`p 20 20 20`p 20 20 R0 R0 20 20 20 20 20 20`p 20 20 �0`pP��  �	
 ��i�  �� �*   b   20 b0`pP      b   b0`pP         b         B0`   B0`   20 20 20 20       20`p b0`                  B   B                                                                                    B         20    B   B            0`p      20`p          20`p    0      20`p                20`p    0      20`p          20`p       B   B0`   20`p B0`pP   B                              20	 b0`
p	P����   20    B0`   20 20 B0`   B0`   B0`   20 B0`      20 B0`   B0`  
 
20`pP� b   R0 b   b0`   B      b   B0`pP   b0`   20 B   B0`   B0`     
 
R0`pP�    B   20`p    B   20`p 20 20    R0 R0 20 20 R0 R0          B0`   r0 B  �	
 ��"-       B0`pP      B0`pP   B0`pP      B0`   B0`     
 
20`pP� 20 B      20`p 20`p    R0 R0 b0`     
 
R0`pP��	
 ��*  X� �     b0`pP  �	
 ��  K!x �      b0`  �	
 ��-O H$   B0`pP   20 20 B0`pP         20 20 R0 R0 20 20 20 20 20 B0`pP   20 20 r
0	`pP���	
 ��k�  �� �*   b   20 b0`pP      b   b0`pP         b         B0`   B0`   20 20 20 20             20�	
 ��  20�	
 ��  20�	
 ��  20 20�	
 ��  20�	
 ��  20 20 ) 0`pP
 
$ 0`p   B0`  �	
 ��9 U   20 B0`pP  �	
 ��  g� �              p   p   B0`pP   B0`pP      20 B0`pP  �	
 ��   i� �           20`p    20`p B0`pP  	 B0`
p	P����   B0`pP   B0`pP      0   20 B0`pP��   20`p                                                                      20 20 20 20 20 20 20 20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��        20�	
 ��  20�	
 ��  20�	
 �� 	 �0`
p	P����  �	
 ��/  N� �     20 B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`  	 �0`
p	P����  �	
 ��-"P� p� ������� �           R
0	`pP��� b0`   B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   B0`            B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   B0`            b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �      b0`pP  �	
 ��0� �� �         b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �            �0 �0          �0 �0   
  0`
p	P����	
 ��e\N  �I� ��� �� �� �����  �� �� �C� �� �� �  �� �        
  0`
p	P����	
 ��qhN  �I� ��� �� �� �����  �� �� �G� �� �� �� �� �  �� �        �x
  0`
p	����P  �	
 ��d�� �d� �      r0 B0`  �	
 ��(5 C   B0`  �	
 ��(5 C   B0`  �	
 ��$1 ?   B0`  �	
 ��$1 ?   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �                     �0 �0 �0 �0 �0   	 �0`
p	P����  
  0`
p	P����
�      �0`
p	����P
 # 0`
p	P����
 - 0`
p	P����                B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <         R0    20�	
 ��        B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �           20�	
 ��     B0`pP  �	
 ��  h� �     B0`pP  �	
 ��  h� �     B0`  �	
 ��. <   B0`  �	
 ��. <   20 20    20    20�	
 �� 
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �   20�	
 ��  20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 B0`pP  �	
 ��%E����  �� �          20`p
��0`
p	����P
 ) 0`
p	P����	 �0`
p	P����  	 �0`
p	P����  
  0`
p	P      ����
  0`
p	P����
  0`
p	P����
  0`
p	P����	
 ��=3G  �� ��� �����  �S� �� �F         
  0`
p	P����	
 ��=3G  �� ��� �����  �S� �� �F           0`pP�а	
 ����� �   x	  0`
p	P����	
 ��D  ��� �  
  0`
p	P����	
 ��HN�  �	� �W  ��� �z  �� �  �D� �  �?� �  �� �  
  0`
p	P����	
 ��?K�  �
�� �  ��� ��  �<� �  �?� �  �� �   
  0`
p	P����	
 ��?K�  �
�� �  ��� ��  �<� �  �?� �  �� �   
  0`
p	P����	
 ��?K�  �
�� �  ��� ��  �<� �  �?� �  �� �   
  0`
p	P����	
 ��HR�  �
� �W  ��� �|  �� �  �E� �  �@� �  �� �  
  0`
p	P����	
 ��HO�  �
� �W  ��� �z  �� �  �E� �  �@� �  �� �            b   �0 �0 �0 �0 �0   	 	 0`  	      0`pP�а	
 ���� �� �� �    �0    b   b   �0 �0 �0 �0 �0     0   h ! 0`pP�	
 ���� �� �� �    �0    b   �0`  �	
 ��(,y ty �      �0`  �	
 ��L,� �� �   �0`  �	
 ��(-z uz �      �0`  �	
 ��L-� �� �  	 x
  0`pP�  �	
 ��
]_� �    	 x
  0`pP�  �	
 ��
]^� �     20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20�	
 ��  20 20 20 20 20 20�	
 ��  20 20 20 20 20 20 20�	
 ��  20�	
 �� 
 
r0`pP��	
 ��$B  a� �  �� �  �� �   �0`pP��  �	
 ��0D  e� �  �� �  �� �  �� ��        �0`  �	
 ��  .!u �      �0`  �	
 ��  ."v �     
 
r0`pP��	
 ��/S  r� �  �� �  �� �  �� �;   
 
r0
      `pP��	
 ��/S  r� �  �� �  �� �  �� �;    �0`pP��  �	
 ��AU  v� �  �� �  �� �  �� �=  �� �� ��     �0`pP��  �	
 ��AU  v� �  �� �  �� �  �� �=  �� �� ��     �0`  �	
 ��$  :_ x   �0`  �	
 ��$  :_ x  
 
�0`pP��	
 ��?  i� x!� �   
 
�0`pP��	
 ��@  j� y"� �                �0 �0  0`pP�  �	
 ��|  ��� �   h
 
 0`p  �	
 ��  ��� �  	 x  0`pP�  �	
 ��x  �� �0   	 x  0`pP�  �	
 ��y  �� �0    20`p�	
 ����  �� �h  �� �� �?  �� �  �� ��  �� �� ��  �	� �	� �
  �
� �
i  �� �� ��  �� �� ��  �� �� ��                                                                           20 20 20 20 20 20 20 20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��        20�	
 ��  20�	
 ��  20�	
 ��  20�	
 �� 	 �0`
p	P����  �	
 ��/  N� �     20 B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`   B0`  	 �0`
p	P����  �	
 ��9/T� �� ������� ���  ��         B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   B0`            B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   B0`            b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �      b0`pP  �	
 ��0� �� �         b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �            �0 �0          �0 �0   
  0`
p	P����	
 ��qhQ{  �Q� ��� �� �� �����  �9� �$� �� �� �� �� �� �  �� �        
  0`
p	P����	
 ��qhQ{  �Q� ��� �� �� �����  �9� �$� �� �� �� �� �� �  �� �        �x
  0`
p	����P  �	
 ��d�� �q� �      r0 B0`  �	
 ��(5 C   B0`  �	
 ��(5 C   B0`  �	
 ��$1 ?   B0`  �	
 ��$1 ?   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         B0`   B0`   B0`   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �                     �0 �0 �0 �0 �0   	 �0`
p	P����  	  
0	`pP      ���  
��0`
p	����P	 $ 
0	`pP���  	 . 
0	`pP���                  B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <         R0    20�	
 ��        B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �           20�	
 ��     B0`pP  �	
 ��  h� �     B0`pP  �	
 ��  h� �     B0`  �	
 ��. <   B0`  �	
 ��. <   20 20    20    20�	
 �� 
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �   20�	
 ��  20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 B0`pP  �	
 ��%E����  �� �          20`p
��0`
p	����P
 ) 0`
p	P����	  
0	`pP���  	  
0	`pP���  
        0`
p	P���� x  0`
p	P����
  0`
p	P����	
 ��A8G  �� ��� �����  �u� �  �� �        
  0`
p	P����	
 ��A8G  �� ��� �����  �u� �  �� �         h 
 0`p  �	
 ����� �   x h
  0`pP�а	
 ��K  ��� �  
  0`
p	P����	
 ��4F�  ��� ��  �#� �  ��� �  �� �2  
  0`
p	P����	
 ��3K�  �
�	� ��  �� �  �9� �  �� �2   
  0`
p	P����	
 ��3K�  ��� ��  �#� �  �q� �  �� �2   
  0`
p	P����	
 ��3K�  �
�� ��  �� �  �8� �  �� �2   
  0`
p	P����	
 ��3R�	  ��	� ��  �� �  �7� �  �� �2   
  0`
p	P����	
 ��3O�	  ��	� ��  �� �  �7� �  �� �2   
  0`
p	P����       20    20 20 20 20       B   b0`   b0`   20 B0`pP   20 20 B   B0`pP            B0`   �0`   �0`   20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20 20
 
20`pP��	
 ��  Z� �    
 
20`pP��	
 ��  Z� �    
 
20`pP��	
 ��  2-� �    
 
20`pP��	
 ��  2-� �     20�	
 ��           B0`   B0`   B0`  �	
 ��  B0`  �	
 ��  B0`  �	
 �� 
 
R0`pP�    20 20
 
20`pP��	
 ��  Z� �    
 
20`pP��	
 ��  Z� �    
 
20`pP��	
 ��  2-� �    
 
20`pP��	
 ��  2-� �     20�	
 ��           B0`   B0`   B0`  �	
 ��  B0`  �	
 ��  B0`  �	
 �� 
 
R0`pP�    20`p 20`p B0`pP   B0`pP   B   B   20 r0`p r0`p �0`pP��   �0`pP��   b0`pP   b0`pP  
 
20`pP�
 
20`pP�      
 
20`pP��	
 ���� �   
 
20`pP��	
 ���� �    B0      `   B0`  
 
R0`pP�    20 20
��0`
p	����P b0`  
  0`
p	P���� b0`pP   �0`   �
0	`pP��� �0`pP   r0`p   
 
20`pP��	
 ��T  �� �   
 
20`pP��	
 ���� �� �      B0`pP  �	
 ��          
 
20`pP��	
 ��G  �� �   
 
20`pP��	
 ���� �� �      B0`pP  �	
 ��          
 
20`pP��	
 ��T  �� �   
 
20`pP��	
 ���� �� �      B0`pP  �	
 ��                
 
20`pP��	
 ���� �   
 
20`pP��	
 ���� �    B0`   B0`  
 
R0`pP�       20
��0`
p	����P b0`  
  0`
p	P���� b0`pP   �0`   �
0	`pP��� �0`pP   r0`p   
 
20`pP��	
 ��T  �� �   
 
20`pP��	
 ���� �� �      B0`pP  �	
 ��          
 
20`pP��	
 ��G  �� �   
 
20`pP��	
 ����       �� �      B0`pP  �	
 ��          
 
20`pP��	
 ��T  �� �   
 
20`pP��	
 ���� �� �      B0`pP  �	
 ��           20 R0`p�	
 ��)(��  �
� �� �   }    ���� 20�	
 ��  20�	
 ��  B0`pP  �	
 ��6  Pq b� �    
 
20`pP��	
 ��~� �� �� �     B0`pP  �	
 ��)  Cd U z  
 
20`pP��	
 ��v� �� �� �     B0`pP  �	
 ��2  Q� �� �� �     B0`pP��  �	
 ���� �� �� �� �      B0`   B0`pP  �	
 ���      B0`pP  �	
 ���      B0`pP  �	
 ���      �0`pP      20 20 20 20 20 20 2
0	`pP���	
 ���� �� �� �N� �     
 
20`pP��	
 ��:  Y� �� �@� �     2
0	`pP���	
 ���� �� �� �N� �     
 
20`pP��	
 ��:  Y� �� �A� �    
 
20`pP��	
 ��1  K� ]N� �   
 
20      `pP��	
 ��>  X� jD� �    B0`pP��  �	
 ���� �� �I� �    B0`pP��  �	
 ��~� �� �F� �    
 
20`pP��	
 ��1  K� ]N� �   
 
20`pP��	
 ��>  X� jE� �    B0`pP��  �	
 ��~� �� �Q� �     B0`pP��  �	
 ���� �� �I� �    20 20 20 B0`  �	
 ��  B0`  �	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  B0`  �	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  B0`  �	
 ��  20�	
 ��  20�	
 ��  20 R0`p�	
 ��)(��  �
� �� �   }    ��� 20�	
 ��  20�	
 ��  B0`pP  �	
 ��6  Pq b� �    
 
20`pP��	
 ���� �� �� �    B0`pP  �	
 ��)  Cd U z  
 
20`pP��	
 ��}� �� �� �     B0`pP  �	
 ��2  Q� �� �� �     B0`pP��  �	
       ���� �� �� �� �      B0`   B0`pP  �	
 ���      B0`pP  �	
 ���      B0`pP  �	
 ���      �0`pP      20 20 20 20 20 20 2
0	`pP���	
 ���� �� �� �G� �     
 
20`pP��	
 ��:  Y� �� �@� �     2
0	`pP���	
 ���� �� �� �G� �     
 
20`pP��	
 ��:  Y� �� �A� �    
 
20`pP��	
 ��1  K� ]N� �   
 
20`pP��	
 ��>  X� jD� �    B0`pP��  �	
 ���� �� �J� �    B0`pP��  �	
 ���� �� �F� �   
 
20`pP��	
 ��1  K� ]N� �   
 
20`pP��	
 ��>  X� jE� �    B0`pP��  �	
 ���� �� �J� �    B0`pP��  �	
 ���� �� �G� �    20 20 20 B0`  �	
 ��  B0`  �	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��        B0`  �	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  B0`  �	
 ��  B   B   B   B   B0`  �	
 ��7 2   B0`  �	
 ��7 2   B0`  �	
 ��7 2   B0`  �	
 ��7 2   B0`  �	
 ��7 2  

R0`P  �	
 ��J  b} x   B0`  �	
 ��7 2   B0`  �	
 ��7 2   B0`  �	
 ��7 2   B0`  �	
 ��7 2         20 20          B      B                                 B   B0`   20`p 20`p B0`   20 20    B0`  
 
R0`pP�
 
R0`pP��	
 ��@� i� �    B0`   B0`  �	
 ��an |   B0`  �	
 ��an |   B0`   B0`  �	
 ��  B0`            B      B                                 B   20 B0`   B   B   20 20    B0`  
 
R0`pP�
 
R0`pP��	
 ��@� i� �    B0      `   B0`  �	
 ��	hu �      B0`  �	
 ��	hu �      B0`   B0`  �	
 ��  B0`         20`p
 
R0`pP� 20`p�	
 ��19@I                B0`   20 20 �0`pP   r0`p    20    20             20 20 20 20    20`p�	
 ��5  U| �      B0`pP  �	
 ��z� �� �      B0`  �	
 ��0  Ou �      20`p�	
 ��u� �� �  
 
20`pP� B0`pP  �	
 ���� �    B0`pP  �	
 ��  B0`pP  �	
 ��     20`p�	
 ��5  U| �      B0`pP  �	
 ���� �� �         B0`  �	
 ��0  Ou �      20`p�	
 ��|� �� �  
 
20`pP� B0`pP  �	
 ���� �    B0`pP  �	
 ��  B0`pP  �	
 ��     20    20       20 20    20`p�	
 ��
y� �           20 20    R0`p    20`p�	
 ��
u� �     20`p       B0`pP  �	
 ���� �    B0`pP  �	
 ��  B0`pP  �	
 ��  B0`pP  �	
 ��5'<���x  �y��
� �  �� �   }    p��� B0`pP  �	
 ��5'<���x  �y��
� �  �� �   }    $���	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       |��� b0`  �	
 ��1#  A�|c  �
� �  �� �   }    8��� R0�	
 ��5$  c��7  �
� �  �� �   }       ���� b0`  �	
 ��5&"*  ���� �� �� �
  �   }     ����
 
R0`pP��	
 ��5&,6  ����  �
� �  �� �   }     `��� R0`p b0`pP  �	
 ��5''�  �7��� �� �� �
  �   }    ��� 20`p R0�	
 ��9)  c�{  �� �� �� �
  �   }      ���� r0�	
 ��1"  Szo/  �
� �  �� �   }     t��� R0`p�	
 ��1#&  J�q7  �
� �  �� �   }    0��� R0`p�	
 ��=-&  o      �  ��  �
� �  �� �   }      ���� b0`  �	
 ��9+#  ���  �� �� �� �
  �   }    ���� R0�	
 ��9*   {��  �� �� �� �
  �   }     L��� r0�	
 ��1"  9Ih(  �
� �  �� �   }     ��� �0`  �	
 ��1#%  a}�  �
� �  �� �   }    ����
 
x �0�	
 ��5$!  o��.  �
� �  �� �   }       ���� �0`p�	
 ��5$   l��.  �
� �  �� �   }       8���    R0`p�	
 ��
+� �^     b0`  �	
 ��9)  V�n  �� �� �� �
  �   }      ����             B0`pP                 	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       @���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       8���   	 	 0`�	
 ��A0        ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       0���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       (���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       п��       20`p�	
 ���� �          20 20    20`p    20`p�	
 ��
|� �     20`p B0`pP  �	
 ���� �    B0`pP  �	
 ��  B0`pP  �	
 ��  B0`pP  �	
 ��5'<���v  �&��
� �  �� �   }    ���� B0`pP  �	
 ��5'<���v  �&��
� �  �� �   }    d���	 	 0`�	
 ��A0  ���  ���  �
� �  ��       �   }       ���	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ���� b0`  �	
 ��1#  A�|c  �
� �  �� �   }    x��� R0�	
 ��1!�  ���
� �  �� �   }      8��� b0`  �	
 ��5&"*  ���� �� �� �
  �   }     ���
 
R0`pP��	
 ��5&,  ����8  �
� �  �� �   }     ���� 20`p
 
R0`pP��	
 ��A1,  ���  �#��� �� �� �
  �   }      @��� B0`   R0�	
 ��9*  h��  �� �� �� �
  �   }     ��� r0�	
 ��-|  �R�
� �  �� �   }    ���� R0`p�	
 ��1#&  J�q7  �
� �  �� �   }    l��� R0`p�	
 ��9+&  ���,  ���
� �  �� �   }     ��� b0`  �	
 ��5&#u  ���� �� �� �
  �   }     غ�� R0�	
 ��5& u  ���� �� �� �
  �   }     ���� r0�	
 ��1"  9Ih(  �
� �  �� �   }     T��� �0`  �	
 ��1#%  a}�  �
�       �  �� �   }    ���
 
x �0�	
 ��5$!  o��.  �
� �  �� �   }       ȹ�� �0`p�	
 ��5$   l��.  �
� �  �� �   }       ����    R0`p�	
 ��
+� �`     b0`  �	
 ��9*  c��  �� �� �� �
  �   }     ��� R
0	`pP���	
 ��QA  f����  �3����� �� �  �  �� �   } }    ���� 20`p               	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       0���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ط��   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       (���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ж��   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       x���   	 	 0`�	
 ��A0  ���  ���  �
� �  ��       �   }        ���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ȵ��   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       p���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ���   	 	 0`�	
 ��A0  ���  ���  �
� �  �� �   }       ����                                                                                        20 20 20 20 20 20 20 20 20 20 20 20 R0 R0 R0 R0 R0 R0 R0 R0 R0 R0 R0 20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  B0`  �	
 ��  20    20 20 B0`  	 �0`
p	P����  �	
 ��5+0  D� a� �������  ��        	 �0`
p	P����  �	
 ��,  E� �           20             20 B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         R0 R0 R0 R0          B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         R0 R0 R0 R0          b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �      b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �            �0 �0          �0 �0          20 B0`  �	
 ��(5 C   B0`  �	
 ��(5 C   B0`  �	
 ��$1 ?   B0`  �	
 ��$1 ?   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A               R0 R0 R0 b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �            �0 �0 �0 �0 �0          r0 r0 �0 r0    B0`  �	
 ��4A O   B0`  �	
 ��4A O   B0`  �	
 ��0= K   B0`  �	
 ��0= K  
 
20`pP��	
 ��Q�q� �  ��      
 
20`pP��	
 ��Q�q� �  ��                                  B0`  �	
 ��                 �0                            �0 �0 �0 �0 �0                   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <         R0    20�	
 ��     R0 B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �           20�	
 ��     B0`pP  �	
 ��  g� �     B0`pP        �	
 ��  g� �     B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �        B0`  �	
 ��. <   B0`  �	
 ��. <   20 20    20    20�	
 �� 
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �   20�	
 ��  20
  0`
p	P����	 �0`
p	P����  
  0`
p	P���� 20 20 20 �
0	`pP���	
 ��ma  K�]�r�������������������������� �    }       20 20 20	 �0`
p	P����  �	
 ����  ������	����������	��	��	��	�i�	���  ��	����	��	��	�� �    }      20	 �0`
p	P����  �	
 ����  ������	����������	��	��	��	�i�	���  ��	����	��	��	�� �    }      20       20 20
  0`
p	P���� 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 0`pP b0`pP   b0`  
  0`
p	P����	
 ��]RE�  ��� ��� �	 � �	� �
����  �� �� �\� �  �� �          
  0`
p	P����	
 ��]RE�  ��� ��� �	 � �	� �
����  �� �� �\� �  �� �          �x	  0`
p	����P  �	
 ��a�� ��� �     r0	 B0`
p	P����   b0`   0   0   B0`pP  �	
 ��%E����  �� �          B0`pP  �	
 ��%E����  �� �         
��0`
p	����P r0 r0� 0`
p	����P  
��0`
p	����P r0 r0
��0`
p	����P r0 r0
��0`
p	����P r0 �0`pP   r0�h  0`
p	����P   �0� 0`
p	����P   �0
��0`
p	����P
��0`
p	���       �P
 # 0`
p	P����
 - 0`
p	P����
 ) 0`
p	P����	 �0`
p	P����  	 �0`
p	P����  
  0`
p	P����
  0`
p	P����	 �0`
p	P����  �	
 ��EA  ��� �
�  �� �  
  0`
p	P����	
 ��6  S�� �   
  0`
p	P����	
 ��6  S�� �     0`pP�  �	
 ��A  ^�� �   
  0`
p	P����	
 ��4F�  �� �(  �	c� �  ��� �  ��� ��   �0 �0
  0`
p	P����
  0`
p	P����	
 ��*F�  �� ��  �	�� �
  ��� ��     �0 �0
  0`
p	P����	
 ��*F�  �� ��  �	�� �
  ��� ��     �0 �0
  0`
p	P����	
 ��*F�  �� ��  �	�� �
  ��� ��     �0 �0
  0`
p	P����	
 ��4I�  �� �(  �
�� �W  ��� �  �� ��   �0 �0
  0`
p	P����	
 ��3I�  �� �  �	� �
G  ��� �  �� ��    �0  0`pP �0
  0`
p	P����	
 !      ��DU  �� ��� �    
  0`
p	P����	
 ��DU  �� ��� �     x  
0	`pP���  �	
 ��G  ��� �   x  0`
p	P����	
 ��D  ��� �  
  0`
p	P����       20    20       20 20    20`p�	
 ��	q �            20 20 B0`   20�	
 ��-N@5  �
� �  �� �   }     ��� �0`  �	
 ��-Jf�  �
� �  �� �   }    ���� r0�	
 ��-C~p5  �
� �  �� �   }     l��� r0�	
 ��-8n`5  �
� �  �� �   }     0���    20`p�	
 ��	m{ �         20 B0`   20`p�	
 ���� �    20`p�	
 ��  B0`  �	
 ��  R0 R0 B0`  �	
 ��  B0`  �	
 ��  r0`p�	
 ��=,  B��� �  �� �� �� ��  }       $��� R0`p�	
 ��=-  ���� �  �� �� �� ��  }      Ԛ�� b0`pP  �	
 ��=,  @����� �� �� �  ��  }       ����   "       B0`         B0`pP                 	 �0`
p	P����  �	
 ��E5$  ���������� �� �� �  ��  }      ���� B   b   b   B0`   B0`   B0`   �0`pP��  �	
 ��I9  ���� �/��
��� �  �� �� ��  }      @���          �0`pP��  �	
 ��I9  ���� �/��
��� �  �� �� ��  }      И��          �0`pP��  �	
 ��I9  ���� �)��
��� �  �� �� ��  }      `���    �0`pP��  �	
 ��I9  ���� �/��
��� �  �� �� ��  }      ����    �0`pP��  �	
 ��I9  ���� �/��
��� �  �� �� ��  }      ����    h 
�0`pP��	
 ��I9!  ���� �/��
��� �  �� �� ��  }      (���      
 
�0`pP��	
 ��I9  ���� �/��
��� �  �� �� ��  }      ���� b   �0`pP��  �	
 ��I9  ���� �/��#      
��� �  �� �� ��  }      T���       20`p�	
 ��
x� �           20 20 B0`   20�	
 ��-N@5  �
� �  �� �   }     ̕�� �0`  �	
 ��-Jf�  �
� �  �� �   }    ���� r0�	
 ��-C~p5  �
� �  �� �   }     P��� r0�	
 ��-8n`5  �
� �  �� �   }     ���    20`p�	
 ��
t� �        20 B0`   20`p�	
 ���� �    20`p�	
 ��  B0`  �	
 ��  R0 R0 B0`  �	
 ��  B0`  �	
 ��  r0`p�	
 ��=,  B��� �  �� �� �� ��  }       ��� b0`pP  �	
 ��=-  �� ���� �  �� �� ��  }      ���� b0`pP  �	
 ��=,  @����� �� �� �  ��  }       `���    20       20`p               	 �0`
p	P����  �	
 ��E4$  �$�����I��� �� �� �  ��  }       Ȓ�� B   B0`   R0 B0`pP��  �	
 ��I8@�$      ���  ���� ���� �� �
  �   } }     H���
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      ���         
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      |���         
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      ���   
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      ����   
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      H���    h �0`pP  �	
 ��I9  ���� ���
��� �  �� �� ��  }      ����        0`pP�	
 ��I9  ���� ���
��� �  �� �� ��  }      x��� b  
 
�0`pP��	
 ��I9  ���� ���
��� �  �� �� ��  }      ���   � 0`
p	����P  2	0`p�P  
 
20`pP�                                          %                         20 20 B0`pP��   2
0	`pP��� 20 20 B0`pP��   2
0	`pP���    B0`pP  �	
 ��VZ h   20    b   b         20 20                                                       20             20 R0`p b      B0`pP  �	
 ��VZ h   20    b   b         20 20                                                       20             20 R0`p b                           B         B0`            B   B                                
 
R0`pP�	 b0`
p	P����   B0`                                       20 20�	
 ��                                                  B0`pP   B  �	
 ��"7                   B   B               b0`pP   b0`pP   20 20&      �	
 ��  20 B0`   B0`     
 
R0`pP� b   b      b   R0 b   b0`   B      b0`  	 b0`
p	P����   b   b   R0 b   b0`   B   b0`   b   b   b   b   B   B   B   b   B   B0`   B   B   b   b0`pP   R0`p b0`pP   b0`         B   B   B0`   B0`   B   B   20             2
0	`pP���    20`p B0`   B0`pP      20`p   
 
20`pP�    20`p    B0`pP      20`p   
 
20`pP�    20`p    B0`pP      20`p    B0`   B0`   B0`   B0`pP  
 
20`pP� B0`              
 
20`pP��	
 ��
;O� �     b0`pP  �	
 ��+1h {   R0`p       R0`p       R0`p       20`p�	
 ��$  3C V         R0`p B   B   B   B  '       B   B         B0`   B0`               20                                                                                           20 20 20 20 20 20 20 20 20 20 20 20 R0 R0 R0 R0 R0 R0 R0 R0 R0 R0 R0 20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  20�	
 ��  B0`  �	
 ��  20    20 20	 �0`
p	P����  �	
 ��A70  E� t� �������  �� ����        	 �0`
p	P����  �	
 ��,  E� �           20       20 B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         R0 R0 R0 R0          B0`  �	
 ��+8 F   B0`  �	
 ��+8 F   B0`  (      �	
 ��'4 B   B0`  �	
 ��'4 B   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         R0 R0 R0 R0          b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �      b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �   b0`pP  �	
 ��0� �� �            �0 �0          �0 �0          20 B0`  �	
 ��(5 C   B0`  �	
 ��(5 C   B0`  �	
 ��$1 ?   B0`  �	
 ��$1 ?   B0`  �	
 ��&3 A   B0`  �	
 ��&3 A         R0 R0 R0 b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �   b0`pP  �	
 ��-� �� �            �0 �0 �0 �0 �0          r0 r0 �0 r0    )      B0`  �	
 ��4A O   B0`  �	
 ��4A O   B0`  �	
 ��0= K   B0`  �	
 ��0= K  
 
20`pP��	
 ��Q�q� �  ��      
 
20`pP��	
 ��Q�q� �  ��                                  B0`  �	
 ��                 �0                            �0 �0 �0 �0 �0                   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <   B0`  �	
 ��. <         R0    20�	
 ��     R0 B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �           20�	
 ��     B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �     B0`pP  �	
 ��  g� �        B0`  �	
 ��. <   B0`  �	
 ��. <   20 20    20    20�	
 �� 
 
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �  
 *      
20`pP��	
 ��%� �� �  
 
20`pP��	
 ��%� �� �   20�	
 ��  20
  0`
p	P����	 �0`
p	P����  	  
0	`pP���   20 20 20 �
0	`pP���	
 ��qg  K�]�r������������������������ �  ����  }     20 20 20	 �0`
p	P����  �	
 ����  ��
��
��	��
��	��
��
��
��
��
��	�k��"  ��
����
����
����	 �	  �	�	�	�	�
�
  }        20	 �0`
p	P����  �	
 ����  ��
��
��	��
��	��
��
��
��
��
��	�k��"  ��
����
����
����	 �	  �	�	�	�	�
�
  }        20 20 20	 ( 
0	`pP���   20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 0`pP�   b0`pP   b0`  
  0`
p	P����	
 ��]RF�  ���+       ��� �	"� �	� �
����  �� �� �h� �  �� �          
  0`
p	P����	
 ��]RF�  ��� ��� �	"� �	� �
����  �� �� �h� �  �� �          �x	  0`
p	����P  �	
 ��`�� �|� �      r0 R
0	`pP��� b0`   0   0   B0`pP  �	
 ��%E����  �� �          B0`pP  �	
 ��%E����  �� �         
��0`
p	����P r0 r0� 0`
p	����P  
��0`
p	����P r0 r0
��0`
p	����P r0 r0
��0`
p	����P r0 �0`pP   r0�h  0`
p	����P   �0� 0`
p	����P   �0
��0`
p	����P
��0`
p	����P	 $ 
0	`pP���  	 . 
0	`pP���  
 ) 0`
p	P����	  
0	`pP���  	  
0	`pP���  
  0`
p	P���� x
  0`
p	P����
  0`
p	P����	
 ��HN  ��	� ��  �� �  
  0`
p	P,      ����	
 ��A  ^�� �   
  0`
p	P����	
 ��A  ^�� �   
  0`
p	P����	
 ��A  ^�� �   
  0`
p	P����	
 ��F�  �� ��  �
�� ��     �0 �0
  0`
p	P����
  0`
p	P����	
 ��F�  �� ��  �
�� ��     �0 �0
  0`
p	P����	
 ��F�  �� ��  �
�� ��     �0 �0
  0`
p	P����	
 ��F�  �� ��  �
�� ��     �0 �0
  0`
p	P����	
 ��I�  �� ��  ��� ��     �0 �0
  0`
p	P����	
 ��I�  �� ��  �
�� ��     �0
 
 0`p   �0
  0`
p	P����	
 ��DU  �� ��� �    
  0`
p	P����	
 ��DU  �� ��� �    	 x	  0`pP�  �	
 ��I  ��� �  ! !x
 h	  
0	`pP���  �	
 ��U  ��� �  
  0`
p	P����                            B         20`p          B   B                             -         
 
R0`pP�	 b0`
p	P����   B0`                                       20 20�	
 ��                                                  B0`pP   B  �	
 ��"7                   B   B               b0`pP   b0`pP   20 20�	
 ��  20 B0`   B0`      b0`pP��   b   b      b   R0 b   b0`   B      b0`  	 �0`
p	P����   b   b   R0 b   b0`   B   b0`   b   b   b   b   B   B0`   B   B   B   b   b   B   B   R0`p b0`pP   b0`pP   b0`         B   B   B0`   B0`   B   B   20             0`p      20`p          20`p    0` 0` 20`p          20`p    0   0   20`p          20`p       B   20 20`p.       B0`pP   B              
 
20`pP��	
 ��
=O� �     b0`pP  �	
 ��-0i |   R0`p       R0`p       R0`p       20`p�	
 ��%  4D W         R0`p B   B   B   B   B   B         R0 R0             20             20       20       20 r0       20 B0`pP   B0`   B0`pP            �0`pP     �	
 ��  20�	
 ��  ����         20�	
 ��  m���          B   B0p  �	
 ��    �	
 ��  2p�	
 ��    �	
 ��  B   B   B   B      20 B   B   B                                             R0`p B   B0`   B0`pP   b   B0`pP  
  0`
p	P����	
 ����  �
��
       
 
�0`pP��	
 ��+0Z4� �  �4�        b   B0`  �	
 ��.     }          B   B   B     /                20 20 20`p 20                   20 20 B  �	
 ��  B   B0`pP��  �	
 ��>  }*� �� �   B0`  �	
 ��!�>������    }     B0`  �	
 ��!�A������    }           20       B   B      20 R0`p	 B0`
p	P����   B0`pP               B         20 R
0	`pP���	 �0`
p	P����  
  0`
p	P���� R0`p�	
 ��)Mk  ���c  �B� �   }     �d��   
 
20`pP�    B0`pP   B0`  �	
 ��5_h         20    B  �	
 ��            20   
 
20`pP� B0`   B0`pP   B0`  �	
 ��&/            �0`   b0`pP��  �	
 ��
0�\�           b0`pP��  �	
 ��
0�\�           �0`pP��  �	
 ��
0��           B`p                              B0`  �	
 ��8 3  T   B0`  �	
 0      ��8 3  T   B0`  �	
 ��	 *   B0`  �	
 ��	 *   B0`  �	
 ��. J   20 B0`  �	
 ��. J   20	 b0`
p	P����   b0`pP��   B  �	
 ��!         B  �	
 ��         b0`pP��   B      B      B      B      b0`   B0`pP        	 �0`
p	P����  �	
 ��M=5  ���:  �����C��� �� �  �� �   }      <a��	 �0`
p	P����  �	
 ��5'9�  �G��� �� �� �
  �   }    �`��	 �0`
p	P����  �	
 ��QA!  h��  �������� �� �  �  �� �   } }    x`��	 b0`
p	P����  �	
 ��M=5  ���9  �������� �� �  �� �   }      `��	 b0`
p	P����  �	
 ��5'=�  �4��� �� �� �
  �   }    �_��    0      20 20 20 20 B0`   B0`   b   b   b0`   b   B   b0`pP      B   B   B   1      B   B0`   B0`   b   b   b0`   b   B   b0`pP      B   B   B   B   B  �	
 ��               R0             20 20 20 20 20 R0 20    20    20    20 B0`  �	
 ��$ 2   20 20 20 20 B0`  �	
 ��$ 2   20 20 20
 
20`pP�
 
20`pP� 2
0	`pP���	
 ��
5��           20 2
0	`pP���	
 ��
5��           20   �	
 ��  20�	
 ��    �	
 ��  20�	
 ��  b0`  �	
 �� - ;   20 20 20 20 b0`  �	
 �� - ;   20 20 20    R0    b     �	
 ��  20�	
 ��  b   R0�	
 ��  20�	
 ��  R0�	
 ��  W p      B         20    20       20 20`p 20�	
 ��  20�	
 ��  R0`p�	
 ��	82u �      B    0`pP�  �	
 ��3f� �� �� �� �2      � �� �  �� �*     0`pP�а	
 ��9r� �� �� �� �� �� �� �  �� �;       0`pP�а	
 ��"r� �� �� �� �� �l      0`pP�  �	
 ��-p� �� �� �� �� �  �� �      B0`  �	
 ��"/ =   B0`  �	
 ��"/ =   20 20 20 20 20 20 20               �	
 ��  20�	
 ��        20�	
 ��                                20 �0`  �	
 ��  $F _   B0`      R0 r0`p�	
 ��(� 3y t+                  B   B   R
0	`pP���	
 ��5'4�  �3��� �� �� �
  �   }    |X�� R
0	`pP���	
 ��5'4�  � ��� �� �� �
  �   }    ,X��       20       B0`pP   B0`pP   0` 20 20 20 20 20`p B0`   B0`      20       20`p B0`pP   20 B0`pP��   b0`pP   b0`pP      3      �0`pP��  
 
R0`pP� B0`   b0`  	 B0`
p	P����   B0`   20 B0`pP   20`p
  0`
p	P���� b0`   B0`pP��  
 
20`pP� r
0	`pP��� 2
0	`pP��� B0`pP   20`p	 B0`
p	P����  �C 0`
p	����P  
 
r0`pP� B     �
  T	  t  d  4  �   20 B   B0`  �	
 ��:>  }   �U��    R0 20 20`p�	
 ��&=    }        b0`         B   B0`           
 
R0`pP�

�0`P   B   B0`      �     	 � x h �0`            b0`  
 
�0`pP�
�b0`
p	����P B  
 
20`pP� 20 B0`pP   B0`pP   20 20          20`p B   B   B   B   B   B   b   B   B                     b         �0`pP��   2p � 0`pP B        
 � 0`
p	P���� 20`p B  
 4      
20`pP�    r0 �   �   �0`   �0`pP   r
0	`pP��� �0`pP  � 0`
p	����P   R0`p �   R0`p R
0	`pP��� �   20`p    20`p R0`p	 B0`
p	P����   20`p B0`   b      b0`   B0`  	 �0`
p	P����      R0, ,� #x h  0`
p	P���� B0`pP��  
 
20`pP� 0`         
  0`
p	P���� �0`pP��      �0`p    0   �0`pP��     
 
�0`pP� �   20 r
0	`pP��� 20`p B0`   b  R	0`p�P  
 
20`pP� �0`  �B0`p��P 20`p �0`   �0`  
�B0`
p	����P �0`pP��  
  0`
p	P���� 20 20`p   	 b0`
p	P����   h	  0`
p	P����	 b0`
p	P����   0`pP�        	 �0`
p	P����   B0`   20 b0`   20 B0`pP   20 2
05      	`pP���
 
20`pP� 2
0	`pP���    B0`pP   0   20`p    2
0	`pP��� b0`pP      `p          20             B0`pP   20 �0`pP                 
 
20`pP�    20`p B0`   b0`pP  	 b0`
p	P����   b0`pP��   �0`   r0`p
 
�0`pP� �0`pP��    0`pP�         b      R0 B0`   B0`pP  
 
20`pP� R0 B0`      B0`                                                   20`p B     
 
20`pP� 20`p B0`   20 20
 
 0`p   20`p �0`pP   20	 B0`
p	P����   20`p	B0`pP�     �� (� �  (�     b0`pP      b   b0`pP  
 
r0`pP� B0`pP��   20`p B0`pP  	 B0`
p	P����         B   B   B   B         b0`   B   20 6      20 20 B0`   20`p B0`   � 0`pP B0`                                             B0`pP   B0`pP   r
0	`pP��� r0`p R0`p b0`         �0`pP   B0`pP   20`p 20 20`p 20`p    b0`      �0`pP  
 
20`pP� 20 B0`   R0`p B0`pP   B0`pP   B0`pP   B0`pP   R0`p �0`pP��   r
0	`pP���                                                                                                                                                                                                                                                                                                                                                                                                                           <�         $ �� �         � t�                     �     :�     H�     X�     l� 7          ��     ��     ��     ��     ��     ��     �     �     *�     D�     V�     p�     ��     ��     ��     ��     ��     ��     �     �     0�     J�     \�     p�     ��     ��     ��     ��     ��     ��     �     �     "�     2�     L�     `�     t�     ��     ��     ��     ��     ��     ��     ��      �     �     .�     >�     X�     n�     ��             ��     ��     ��     ��     ��     ��      �     �     �     .�     B�     L�     Z�     l�     v�     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��      �     
�     �      �     *�     4�     >�     F�     P�     X�     b�     l�     v�     ~�     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��                       "      ,      6      @      J      R      Z      d      p      z      �      �      �      �      �      �      �      �      �  8          �      �      �                     $     0     :             �     :�     H�     X�     l�     ��     ��     ��     ��     ��     ��     �     �     *�     D�     V�     p�     ��     ��     ��     ��     ��     ��     �     �     0�     J�     \�     p�     ��     ��     ��     ��     ��     ��     �     �     "�     2�     L�     `�     t�     ��     ��     ��     ��     ��     ��     ��      �     �     .�     >�     X�     n�     ��             ��     ��     ��     ��     ��     ��      �     �     �     .�     B�     L�     Z�     l�     v�     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��      �     
�     �      �     *�     4�     >�     F�     P�     X�     b�     l�     v�     ~�     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��                       "      ,      6      @  9          J      R      Z      d      p      z      �      �      �      �      �      �      �      �      �      �      �      �                     $     0     :              AddVectoredExceptionHandler � CloseHandle � CreateEventA  � CreateSemaphoreA  DeleteCriticalSection +DuplicateHandle 1EnterCriticalSection  GetCurrentProcess GetCurrentProcessId GetCurrentThread  GetCurrentThreadId  _GetHandleInformation  bGetLastError  �GetProcessAffinityMask  �GetStartupInfoA �GetSystemTimeAsFileTime �GetThreadContext  GetThreadPriority GetTickCount  `InitializeCriticalSection zIsDBCSLeadByteEx  {IsDebuggerPresent �LeaveCriticalSection  �MultiByteToWideChar OutputDebugStringA  FQueryPerformanceCounter YRaiseException  �ReleaseSemaphore  �RemoveVectoredExceptionHandler  �ResetEvent  �ResumeThread  �RtlAddFunctionTable �RtlCaptureContext �RtlLookupFunctionEntry  �RtlUnwindEx �RtlVirtualUnwind  �SetEvent  SetLastError  SetProcessAffinityMa:      sk  +SetThreadContext  4SetThreadPriority CSetUnhandledExceptionFilter QSleep YSuspendThread `TerminateProcess  rTlsAlloc  tTlsGetValue uTlsSetValue {TryEnterCriticalSection �UnhandledExceptionFilter  �VirtualProtect  �VirtualQuery  �WaitForMultipleObjects  �WaitForSingleObject �WideCharToMultiByte �__C_specific_handler  @ ___lc_codepage_func C ___mb_cur_max_func  P __doserrno  R __getmainargs S __initenv T __iob_func  [ __lconv_init  ^ __pioinfo a __set_app_type  c __setusermatherr  s _acmdln { _amsg_exit  � _beginthreadex  � _cexit  � _endthreadex  � _errno  � _fdopen � _filelengthi64  � _fileno � _fileno � _fmode  _fstat64  K_initterm �_lseeki64 c_onexit �_read �_setjmp �_strdup �_strnicmp $_ultoa  �_write  �_write  abort calloc  'exit  +fclose  .fflush  0fgetpos 8fopen :fprintf <fputc =fputs @fread Afree  Hfsetpos Mfwrite  Pgetc  Qgetchar Ugetwc bisspace hiswctype  ulocaleconv  {longjmp |malloc  �memchr  �memcmp  �memcpy  �memmove �memset  ;      �printf  �putc  �putwc �realloc �setlocale �setvbuf �signal  �sprintf �strcmp  �strcoll �strerror  �strftime  �strlen  �strncmp �strtoul �strxfrm �towlower  �towupper  �ungetc  �ungetwc �vfprintf  �wcscoll �wcsftime  �wcslen  wcsxfrm  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � KERNEL32.dll    � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � msvcrt.dll                                                                                                                          0@                     @     p�@             <              ��@     p�@     ��A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ,             P@     �                       =      ,    c�       @     u                       ,    ��       �@     2                           ��                      ,    ��      `�@     '                      ,    �b      ��@     z                                                                                                                                                                                                                                                                      _�       GNU C++11 8.1.0 -mtune=core2 -march=nocona -g -std=c++11 F:\debug\ClionWork\EFS\OS\main.cpp F:\debug\ClionWork\EFS\cmake-build-debug P@     �           __builtin_va_list �   char �   size_t #,�   long long unsigned int long long int �   intptr_t >#�   uintptr_t K,�   wint_t j<  short unsigned int <  wctype_t k<  int h  long int pthreadlocinfo �(�  �  threadlocaleinfostruct `��  	 �
  
locale ��   
wlocale ��  �   �
�  
wrefcount �
�   �   �h   
lc_codepa>      ge ��  
lc_collate_cp ��  
lc_handle ��  
lc_id ��  $
lc_category ��  Hlc_clike �h  mb_cur_max �h  lconv_intl_refcount ��  lconv_num_refcount ��  lconv_mon_refcount ��   lconv ��  (ctype1_refcount ��  0ctype1 ��  8pctype ��  @pclmap ��  Hpcumap ��  Plc_time_curr ��  X pthreadmbcinfo �%�  �  threadmbcinfostruct localeinfo_struct �  
locinfo ��   
mbcinfo ��   _locale_tstruct ��  tagLC_ID �t  
wLanguage �<   
wCountry �<  
wCodePage �<   LC_ID �%  �   �  �  wchar_t �  h  unsigned int �  �  �    long unsigned int �  t  �  �    �    �    lconv X-
�  decimal_point .�   thousands_sep /�  grouping 0�  int_curr_symbol 1�  currency_symbol 2�   mon_decimal_point 3�  (mon_thousands_sep 4�  0mon_grouping 5�  8positive_sign 6�  @negative_sign 7�  Hint_frac_digits 8
�   Pfrac_di?      gits 9
�   Qp_cs_precedes :
�   Rp_sep_by_space ;
�   Sn_cs_precedes <
�   Tn_sep_by_space =
�   Up_sign_posn >
�   Vn_sign_posn ?
�   W   <  R  �  unsigned char �  __lc_time_data �  std G qn  __cxx11 
A�N  basic_string<char, std::char_traits<char>, std::allocator<char> >  M�N  *  �^  �a   *  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC4EPcRKS3_ �  �  �  ^  ��   *  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC4EPcOS3_ ?  O  �  ^  ��   _M_p �
^    �  \0wu  ��  _M_local_buf �5��  _M_allocated_capacity ��       X2�u  �  npos e�  _M_dataplus �a   _M_string_length ��  k   _M_data �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc R	  ]	  
�  ^    _M_length �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy �	  �	  
�  �   !_M_data �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv ^  
  
 @       �   "=   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv ^  z
  �
  
�   �  ]5�u  "=   �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv �
  �
  �
  �    _M_capacity �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy L  W  
�  �    _M_set_length �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy �  �  
�  �   !_M_is_local �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv %�  %  +  �   !_M_create �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy ^  �  �  
�  �  �    _M_dispose �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv �  �  
�    _M_destroy �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy U  `  
�  �    _M_construct_aux_2 �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc �  �  
�  �  �    #_M_construct _ZNSt7__cxx1112basic_stringIcSt11cA      har_traitsIcESaIcEE12_M_constructEyc =  M  
�  �  �    �  W#_  M  _Char_alloc_type P�u  $d   _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv �  �  �  
�   $d   _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv "�  =  C  �   %_M_check +_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc �  �  �  �  �  
�   #_M_check_length 5_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc   2  �  �  �  
�   %_M_limit >_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy �  �  �  �  �  �   %_M_disjunct F_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc %�      �  
�   &_S_copy O_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy u  �  
�  �   &_S_move X_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy �  �  
�  �   &_S_assign a_ZNSt7__cxx1112basic_stringIcSB      t11char_traitsIcESaIcEE9_S_assignEPcyc C  �  �  �    '  t_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ �  �  �  �   �   ^D�u  '  x_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcS4_EESA_ n  �  n  n      `}}  '  }_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcS5_S5_ �  �  �  �   '  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ Q  �  
�  
�   (_S_compare �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy h  �  �  �   #_M_assign �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_assignERKS4_   !  
�  (�   #_M_mutate �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy   �  
�  �  �  
�  �   #_M_erase �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy �    
�  �  �  C       )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4Ev M  S  
�   *�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS3_ �  �  
�  ��   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_ �  	  
�  (�   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yRKS3_ _  t  
�  (�  �  ��   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yy �  �  
�  (�  �  �   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yyRKS3_ 2  L  
�  (�  �  �  ��   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EPKcyRKS3_ �  �  
�  
�  �  ��   )�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EPKcRKS3_     
�  
�  ��   )�   _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EycRKS3_ j    
�  �  �   ��   )�   _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EOS4_ �  �  
�  .�   )�   ._ZNSt7__cxx1112basic_sD      tringIcSt11char_traitsIcESaIcEEC4ESt16initializer_listIcERKS3_ @  P  
�  g  ��   )�   2_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_RKS3_ �  �  
�  (�  ��   )�   6_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EOS4_RKS3_ 	    
�  .�  ��   +~basic_string �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED4Ei o  z  
�  h   ,o  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSERKS4_ 4�  �  �  
�  (�   ,o  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEPKc 4�  +  6  
�  
�   ,o  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc 4�  �  �  
�  �    ,o  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ 4�  �  �  
�  .�   ,o  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE 4�  U  `  
�  g   -begin '_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv �  �  �  
�   -begin /_ZNKSt7__cxx1112basic_stringIcSt11char_trE      aitsIcESaIcEE5beginEv n      �   -end 7_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv �  k  q  
�   -end ?_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv n  �  �  �   .reverse_iterator b0�h  -rbegin H_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv �  <  B  
�   .const_reverse_iterator a5Ni  -rbegin Q_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv B  �  �  �   -rend Z_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv �        
�   -rend c_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv B  p   v   �   -cbegin l_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv n  �   �   �   -cend t_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv n  *!  0!  �   -crbegin }_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv B  �!  �!  �   -crend �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv B  �!  �!  F      �   -size �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv �  C"  I"  �   ,[  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv �  �"  �"  �   ,�  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8max_sizeEv �  �"  #  �   +resize �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc X#  h#  
�  �  �    +resize �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEy �#  �#  
�  �   +shrink_to_fit �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv *$  0$  
�   -capacity �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv �  �$  �$  �   +reserve �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy �$  �$  
�  �   +clear �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv F%  L%  
�   -empty �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv %�  �%  �%  �   W  [7�u  ,�  _ZNKSt7__cxx1112basic_stringIcSt1G      1char_traitsIcESaIcEEixEy �%  &  &  �  �   B  Z2�u  ,�  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy &  o&  z&  
�  �   -at )_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy �%  �&  �&  �  �   -at >_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy &  &'  1'  
�  �   -front N_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv &  �'  �'  
�   -front Y_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv �%  �'  �'  �   -back d_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv &  >(  D(  
�   -back o_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv �%  �(  �(  �   ,  }_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ 4�  �(  �(  
�  (�   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc 4�  P)  [)  
�  
�   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc 4�  �)  �)  
�  �    ,  �_ZNSt7__cxx1112basic_striH      ngIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE 4�  *  '*  
�  g   ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ 4�  �*  �*  
�  (�   ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy 4�  �*  �*  
�  (�  �  �   ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy 4�  S+  c+  
�  
�  �   ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKc 4�  �+  �+  
�  
�   ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc 4�  ,  +,  
�  �  �    ,�   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendESt16initializer_listIcE 4�  �,  �,  
�  g   +push_back 2_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9push_backEc �,  -  
�  �    ,�  A_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ 4�  _-  j-  
�  (�   ,�  Q_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ 4�  �-  �-  
�  .�   ,�I        h_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy 4�  (.  =.  
�  (�  �  �   ,�  x_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKcy 4�  �.  �.  
�  
�  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc 4�  �.  /  
�  
�   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc 4�  ]/  m/  
�  �  �    ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE 4�  �/  �/  
�  g   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc �  `0  u0  
�  n  �  �    )�  8_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE 1  1  
�  �  g   ,�  L_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ 4�  l1  |1  
�  �  (�   ,�  c_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_J      yy 4�  �1  �1  
�  �  (�  �  �   ,�  z_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy 4�  K2  `2  
�  �  
�  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKc 4�  �2  �2  
�  �  
�   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc 4�  3  43  
�  �  �  �    ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEc �  �3  �3  
�  �3  �    __const_iterator ln  -erase �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy 4�  04  @4  
�  �  �   -erase _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE �  �4  �4  
�  �3   -erase _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ �  F5  V5  
�  �3  �3   +pop_back ,_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv �5  �5  
�   ,   E_ZNK      St7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ 4�  6  %6  
�  �  �  (�   ,   [_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_yy 4�  �6  �6  
�  �  �  (�  �  �   ,   t_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy 4�  �6  7  
�  �  �  
�  �   ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc 4�  q7  �7  
�  �  �  
�   ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc 4�  �7  �7  
�  �  �  �  �    ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ 4�  }8  �8  
�  �3  �3  (�   ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y 4�  9  /9  
�  �3  �3  
�  �   ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ 4�  �9  �9  
�  �L      3  �3  
�   ,   �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc 4�  G:  a:  
�  �3  �3  �  �    ,   /_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ 4�  �:  �:  
�  �3  �3  �  �   ,   :_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ 4�  �;  �;  
�  �3  �3  
�  
�   ,   E_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ 4�  ,<  F<  
�  �3  �3  �  �   ,   P_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ 4�  �<  �<  
�  �3  �3  n  n   ,   i_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE 4�  {=  �=  
�  n  n  g   %_M_replace_aux �_ZNSt7__cxx1M      112basic_stringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc 4�  �=  >  
�  �  �  �  �    %_M_replace �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replaceEyyPKcy 4�  z>  �>  
�  �  �  
�  �   %_M_append �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy 4�  �>  ?  
�  
�  �   -copy �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy �  \?  q?  �  �  �  �   +swap �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ �?  �?  
�  4�   -c_str �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5c_strEv 
�  &@  ,@  �   -data �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv 
�  �@  �@  �   -get_allocator �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv M  �@  �@  �   ,  	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy �  MA  bA  �  
�  �  �   ,  	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERN      KS4_y �  �A  �A  �  (�  �   ,  <	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy �  "B  2B  �  
�  �   ,  M	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy �  �B  �B  �  �   �   ,�  Z	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y �  �B  C  �  (�  �   ,�  |	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy �  ZC  oC  �  
�  �  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy �  �C  �C  �  
�  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy �  -D  =D  �  �   �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y �  �D  �D  �  (�  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcyy �  E  'E  �  
�  �  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy �  �E  �E  �  
�  �   ,�  �	O      _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEcy �  �E  F  �  �   �   ,  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y �  iF  yF  �  (�  �   ,   
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy �  �F  �F  �  
�  �  �   ,  .
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcy �  OG  _G  �  
�  �   ,  B
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy �  �G  �G  �  �   �   ,�  P
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofERKS4_y �  4H  DH  �  (�  �   ,�  s
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy �  �H  �H  �  
�  �  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy �  $I  4I  �  
�  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy �  �I  �I  P      �  �   �   ,�   �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y �  J  J  �  (�  �   ,�   �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy �  �J  �J  �  
�  �  �   ,�   �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy �  �J  K  �  
�  �   ,�   �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEcy �  mK  }K  �  �   �   -substr �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy   �K  �K  �  �  �   ,R   _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ h  BL  ML  �  (�   ,R   e_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ h  �L  �L  �  �  �  (�   ,R   _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy h  M  =M  �  �  �  (�  �  �   ,R   �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEPKc h  �MQ        �M  �  
�   ,R   �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc h  �M  N  �  �  �  
�   ,R   �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKcy h  mN  �N  �  �  �  
�  �   /�  �   0�   JY  0�  �a     string J!   1
A  2@��  2�-  2���  2�҉  2��  2��  2�5�  2�Z�  2�x�  2���  2���  2�Ԋ  2��  2��  2�E�  2�f�  2���  2���  2�ҋ  2��  2��  2�0�  2�P�  2�w�  2���  2���  2��  2��  2�)�  2�I�  2�n�  2���  2���  2�ɍ  2��  2��  2�7�  2�P�  2�t�  2���  2���  2��  2��  2�;�  2�c�  2���  2���  2�ʏ  2��  2��  2�,�  2�Q�  2�w�  2���  2���  2�Ӑ  2��  2��  2�/�  2�M�  3r�  3	��  3
Ƒ  3;�  3w�  3�  3!)�  3%r�  3&��  3'Ƒ  u   V
0Q  4u   Y_ZNSt9nothrow_tC4Ev )Q  �    �P  5nothrow ]_ZSt7nothrow 0Q  6__exception_ptr 	4�U  7�  	O�U  _M_exception_objR      ect 	Q�   8�  	S_ZNSt15__exception_ptr13exception_ptrC4EPv �Q  �Q  ��  �    _M_addref 	U_ZNSt15__exception_ptr13exception_ptr9_M_addrefEv "R  (R  ��    _M_release 	V_ZNSt15__exception_ptr13exception_ptr10_M_releaseEv sR  yR  ��   !_M_get 	X_ZNKSt15__exception_ptr13exception_ptr6_M_getEv �  �R  �R  ��   9�  	`_ZNSt15__exception_ptr13exception_ptrC4Ev S  S  ��   9�  	b_ZNSt15__exception_ptr13exception_ptrC4ERKS0_ FS  QS  ��   �   9�  	e_ZNSt15__exception_ptr13exception_ptrC4EDn �S  �S  ��  EV   9�  	i_ZNSt15__exception_ptr13exception_ptrC4EOS0_ �S  �S  ��  �   :o  	v_ZNSt15__exception_ptr13exception_ptraSERKS0_ �  $T  /T  ��   �   :o  	z_ZNSt15__exception_ptr13exception_ptraSEOS0_ �  qT  |T  ��  �   ;~exception_ptr 	�_ZNSt15__exception_ptr13exception_ptrD4Ev �T  �T  ��  h   ;swap 	�_ZNSt15__exception_ptr13exception_ptr4swapERS0_ U  U  ��  �   <operator bool 	�_ZNKSt15__exception_ptr13exception_ptrcvbEv %�  eU  kU  ��   =__cxa_exception_typeS       	�_ZNKSt15__exception_ptr13exception_ptr20__cxa_exception_typeEv 2�  �U  ��    jQ  2	I�U   2	9jQ  >rethrow_exception 	E_ZSt17rethrow_exceptionNSt15__exception_ptr13exception_ptrE EV  jQ   nullptr_t 
��  ?type_info WV  integral_constant<bool, false> E2W  @value G--�  A�  H-%�  !operator std::integral_constant<bool, false>::value_type J_ZNKSt17integral_constantIbLb0EEcvbEv �V  W  W  8�   B_Tp %�  C__v %�    gV  integral_constant<bool, true> E X  @value G--�  A�  H-%�  !operator std::integral_constant<bool, true>::value_type J_ZNKSt17integral_constantIbLb1EEcvbEv lW  �W  �W  >�   B_Tp %�  C__v %�   7W  D__swappable_details u	__is_integer<long double> `X  E�  �VX  F+     B_Tp ��   __is_integer<double> �X  E�  ��X  F+     B_Tp +�   __is_integer<float> �X  E�  ��X  F+     B_Tp Z�   �   L
Y  4�   L+_ZNSt21piecewise_construct_tC4Ev Y  S�    �X  Gpiecewise_construct O5Y   H__debug 2char_traits<char> �\  '�  _ZNSt11chT      ar_traitsIcE6assignERcRKc �Y  {�  ��   IQ  !�   �Y  (eq  _ZNSt11char_traitsIcE2eqERKcS2_ %�  �Y  ��  ��   (lt $_ZNSt11char_traitsIcE2ltERKcS2_ %�  )Z  ��  ��   JR   ,_ZNSt11char_traitsIcE7compareEPKcS2_y h  pZ  ��  ��  �\   J[  :_ZNSt11char_traitsIcE6lengthEPKc �\  �Z  ��   J  D_ZNSt11char_traitsIcE4findEPKcyRS1_ ��  �Z  ��  �\  ��   (move R_ZNSt11char_traitsIcE4moveEPcPKcy ��  1[  ��  ��  �\   (copy Z_ZNSt11char_traitsIcE4copyEPcPKcy ��  u[  ��  ��  �\   J�  b_ZNSt11char_traitsIcE6assignEPcyc ��  �[  ��  �\  �Y   Jb  j_ZNSt11char_traitsIcE12to_char_typeERKi �Y  �[  ��   Ig  !h  �[  J�  p_ZNSt11char_traitsIcE11to_int_typeERKc �[  G\  ��   J  t_ZNSt11char_traitsIcE11eq_int_typeERKiS2_ %�  �\  ��  ��   Keof x_ZNSt11char_traitsIcE3eofEv �[  (not_eof |_ZNSt11char_traitsIcE7not_eofERKi �[  �\  ��   /�  �    size_t 
��   char_traits<wchar_t> ��`  '�  �_ZNSt11char_traitsIwE6assignERwRKw f]  ��  ��   IQ  �!�U        f]  (eq �_ZNSt11char_traitsIwE2eqERKwS2_ %�  �]  ��  ��   (lt �_ZNSt11char_traitsIwE2ltERKwS2_ %�  �]  ��  ��   JR   �_ZNSt11char_traitsIwE7compareEPKwS2_y h  5^  ��  ��  �\   J[  �_ZNSt11char_traitsIwE6lengthEPKw �\  m^  ��   J  �_ZNSt11char_traitsIwE4findEPKwyRS1_ ��  �^  ��  �\  ��   (move �_ZNSt11char_traitsIwE4moveEPwPKwy ��  �^  ��  ��  �\   (copy �_ZNSt11char_traitsIwE4copyEPwPKwy ��  :_  ��  ��  �\   J�  �_ZNSt11char_traitsIwE6assignEPwyw ��  }_  ��  �\  f]   Jb  �_ZNSt11char_traitsIwE12to_char_typeERKt f]  �_  ��   Ig  �!-  �_  J�  �_ZNSt11char_traitsIwE11to_int_typeERKw �_  `  ��   J  �_ZNSt11char_traitsIwE11eq_int_typeERKtS2_ %�  R`  ��  ��   Keof �_ZNSt11char_traitsIwE3eofEv �_  (not_eof �_ZNSt11char_traitsIwE7not_eofERKt �_  �`  ��   /�  �   20��  21֒  22��  23�  25�  26�  27?�  28j�  2:9�  2;d�  2<��  2=��  2?��  2@
  2Bƒ  2C�  2D�  2E(�  2G��  2H)�  2IT�V        2J�  2LN�  2Mz�  2N��  2Oԓ  2Q��  2R  25  26�  27�  ptrdiff_t 
��   allocator<char> lib  L�n   93   �_ZNSaIcEC4Ev 
b  b  ��   93   �_ZNSaIcEC4ERKS_ 1b  <b  ��  ��   M~allocator �_ZNSaIcED4Ei ]b  ��  h    �a  2Ӗ  2��  2�ݘ  2���  2��  2�'�  2�?�  2���  2���  2���  2�ۙ  2���  2��  2�C�  2�g�  2�u�  2���  2���  2�͚  2��  2��  2�1�  2���  2�*r  2�P�  2�n�  2�қ  2���  2���  2��  2b��  2cД  2e�  2f)�  2gC�  2h[�  2iu�  2j��  2k��  2lΜ  2m�  2n�  2q0�  2rX�  2s}�  2t��  2u��  2v�  2x��  2y�  2|(�  2~@�  2V�  2�q�  2���  2���  2���  2�؞  2��  2��  2�>�  2�^�  2�o�  2���  2���  2�Ο  2��  2��  2�;�  2�`�  2��  2���  allocator_traits<std::allocator<char> > �g  I�  ��  J�  �_ZNSt16allocator_traitsISaIcEE8allocateERS0_y �d  7e  Р  Ie   I�  �,�a  7e  I    �$�\  J�  �_W      ZNSt16allocator_traitsISaIcEE8allocateERS0_yPKv �d  �e  Р  Ie  �e   const_void_pointer �-v�  '(  �_ZNSt16allocator_traitsISaIcEE10deallocateERS0_Pcy f  Р  �d  Ie   J�  �_ZNSt16allocator_traitsISaIcEE8max_sizeERKS0_ Ie  Yf  ֠   (select_on_container_copy_construction �_ZNSt16allocator_traitsISaIcEE37select_on_container_copy_constructionERKS0_ 7e  �f  ֠   I�  ��   I�  �'
�  rebind_alloc �%�a  /�  �a   initializer_list<char> /�h  �   6
�  _M_array :8g       5�\  _M_len ;Wg  �  >_ZNSt16initializer_listIcEC4EPKcy �g  �g  :�  �g  Wg      7
�  9�  B_ZNSt16initializer_listIcEC4Ev �g  �g  :�   Nsize G_ZNKSt16initializer_listIcE4sizeEv Wg  2h  8h  @�   Nbegin K_ZNKSt16initializer_listIcE5beginEv �g  sh  yh  @�   Nend O_ZNKSt16initializer_listIcE3endEv �g  �h  �h  @�   B_E �    g  ?reverse_iterator<__gnu_cxx::__normal_iterator<char*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > > ?reverse_iX      terator<__gnu_cxx::__normal_iterator<char const*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > > O_V2 GPG�i  Qios_base �j  RInit [+Init __ZNSt8ios_base4InitC4Ev 3j  9j  F�   +~Init `_ZNSt8ios_base4InitD4Ev ej  pj  F�  h   S_S_refcount ca�  S_S_synced_with_stdio d%�    2RL�  2SW  2T-  2\^�  2e�  2h��  2i��  Qbasic_ostream<char, std::char_traits<char> > "k  /�  �   0�   JY   Qbasic_ostream<wchar_t, std::char_traits<wchar_t> > mk  /�  �  0�   ]   Qbasic_istream<char, std::char_traits<char> > �k  /�  �   0�   JY   Qbasic_istream<wchar_t, std::char_traits<wchar_t> > �k  /�  �  0�   ]   istream �!mk  5cin <_ZSt3cin �k  ostream �!�j  5cout =_ZSt4cout "l  5cerr >_ZSt4cerr "l  5clog ?_ZSt4clog "l  wistream �#�k  5wcin B_ZSt4wcin wl  wostream �#"k  5wcout C_ZSt5wcout �l  5wcerr D_ZSt5wcerr �l  5wclog E_ZSt5wclog �l  T__ioinit J�i  Uabs N_ZSt3abse ��  ,m  ��   Uabs J_ZSt3absf Z�  Lm  Z�   UabsY       F_ZSt3absd +�  lm  +�   Uabs =_ZSt3absx �   �m  �    Uabs 8_ZSt3absl t  �m  t   Udiv �_ZSt3divll �  �m  t  t   iterator_traits<char*> � n  A�  �+�a  A�  �+�  AB  �+��  /Z   �   Viterator_traits<char const*> �A�  �+�a  A�  �+
�  AB  �+��  /Z   
�    W__gnu_cxx 
��  X__cxx11 
A1
A�n  2�r�  3��  3Ƒ  H__ops #2,�\  2-�a  new_allocator<char> :�q  9y  O_ZN9__gnu_cxx13new_allocatorIcEC4Ev  o  &o  }�   9y  Q_ZN9__gnu_cxx13new_allocatorIcEC4ERKS1_ _o  jo  }�  ��   ;~new_allocator V_ZN9__gnu_cxx13new_allocatorIcED4Ev �o  �o  }�  h   �  ?�  Naddress Y_ZNK9__gnu_cxx13new_allocatorIcE7addressERc �o  p  p  ��  p   B  A��  �  @
�  Naddress ]_ZNK9__gnu_cxx13new_allocatorIcE7addressERKc p  rp  }p  ��  }p   W  B��  :�  c_ZN9__gnu_cxx13new_allocatorIcE8allocateEyPKv �o  �p  �p  }�  �p  v�       =�\  9(  t_ZN9__gnu_cxx13new_allocatorIcE10deallocateEPcy +q  ;q  }�  �o  �p   :�  �_ZNK9Z      __gnu_cxx13new_allocatorIcE8max_sizeEv �p  |q  �q  ��   B_Tp �    �n  __numeric_traits_integer<int> 7�q  Yy  :o  Y$  ;o  Y�   ?-�  Y�  @o  /K   h   2���  2�P�  2�n�  2���  2���  2�қ  2��  Udiv �_ZN9__gnu_cxx3divExx ��  Zr  �   �    2��  2�;�  2�`�  2��  2���  __alloc_traits<std::allocator<char>, char>  2
�u  2 2
Ve  2 2
�d  2 2
�e  2 2
f  �d   U_S_select_on_copy  ^_ZN9__gnu_cxx14__alloc_traitsISaIcEcE17_S_select_on_copyERKS1_ �a  ?s  ��   Z_S_on_swap  a_ZN9__gnu_cxx14__alloc_traitsISaIcEcE10_S_on_swapERS1_S3_ �s  ܠ  ܠ   [_S_propagate_on_copy_assign  d_ZN9__gnu_cxx14__alloc_traitsISaIcEcE27_S_propagate_on_copy_assignEv %�  [_S_propagate_on_move_assign  g_ZN9__gnu_cxx14__alloc_traitsISaIcEcE27_S_propagate_on_move_assignEv %�  [_S_propagate_on_swap  j_ZN9__gnu_cxx14__alloc_traitsISaIcEcE20_S_propagate_on_swapEv %�  [_S_always_equal  m_ZN9__gnu_cxx14__alloc_traitsISaIcEcE15_S_always_equalEv %�  [_S_nothrow_move  p_ZN9__gnu_cxx14__alloc_[      traitsISaIcEcE15_S_nothrow_moveEv %�  A�   :5�f  fu  A�   ;5�d  A�   <5�f  A     =5Ie  AB   @5�  AW   A5�  rebind<char>  t�u  other  uA�f  B_Tp �    /�  �a   \__normal_iterator<char*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > !�x}  ]  !��   )�  !_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4Ev �v  �v  o�   *�  !_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4ERKS1_ Ww  bw  o�  u�   ^B  !2
n  ,3  !_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEdeEv bw  �w  �w  {�   ^�  !2�m  ,�   !_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEptEv �w  lx  rx  {�   ,�  !!_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEv ��  �x  �x  o�   ,�  !(_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11ch\      ar_traitsIcESaIcEEEEppEi �u  ^y  iy  o�  h   ,   !-_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEv ��  �y  �y  o�   ,   !4_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEi �u  Uz  `z  o�  h   ,�  !9_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEixEx bw  �z  �z  {�  �z   ^�  !8�m  ,  !=_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEpLEx ��  `{  k{  o�  �z   ,=  !A_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEplEx �u  �{  �{  {�  �z   ,�   !E_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmIEx ��  ]|  h|  o�  �z   ,G  !I_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmiEx �u  �|  �|  {�  �z   -base !M_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIc]      St11char_traitsIcESaIcEEEE4baseEv u�  _}  e}  {�   /Z   �  /7     �u  \__normal_iterator<char const*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > !��  ]  !�
�   )�  !_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4Ev w~  }~  W�   *�  !_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4ERKS2_ �~  �~  W�  ]�   ^B  !2Zn  ,3  !_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEdeEv �~    �  c�   ^�  !2Nn  ,�   !_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEptEv �  �  �  c�   ,�  !!_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEv i�  ��  ��  W�   ,�  !(_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEi }}  ��  �  W�  h   ,   !-_ZN9__gnu_cxx17__normal_^      iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEv i�  {�  ��  W�   ,   !4_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEi }}  ��   �  W�  h   ,�  !9_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEixEx �~  u�  ��  c�  ��   ^�  !8Bn  ,  !=_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEpLEx i�  �  �  W�  ��   ,=  !A_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEplEx }}  ��  ��  c�  ��   ,�   !E_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmIEx i�  �  �  W�  ��   ,G  !I_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmiEx }}  ��  ��  c�  ��   -base !M_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEE4baseEv ]�  �  �  c�   /Z   
�  /7     }_      }  __numeric_traits_floating<float> d��  Y  go  Y�   j-�  YL  ko  Y�  lo  /K   Z�   __numeric_traits_floating<double> d�  Y  go  Y�   j-�  YL  ko  Y�  lo  /K   +�   __numeric_traits_floating<long double> dV�  Y  go  Y�   j-�  YL  ko  Y�  lo  /K   ��   __numeric_traits_integer<long unsigned int> 7ņ  Yy  :�  Y$  ;�  Y�   ?-�  Y�  @o  /K   �   __numeric_traits_integer<char> 7'�  Yy  :�   Y$  ;�   Y�   ?-�  Y�  @o  /K   �    __numeric_traits_integer<short int> 7��  Yy  :�  Y$  ;�  Y�   ?-�  Y�  @o  /K   ܈   V__numeric_traits_integer<long long int> 7Yy  :  Y$  ;  Y�   ?-�  Y�  @o  /K   �     _iobuf 0")
��  _ptr "*�   _cnt "+	h  _base ",�  _flag "-	h  _file ".	h  _charbuf "/	h   _bufsiz "0	h  $_tmpfname "1�  ( FILE "3��  ___imp__pctype "���  �  ___imp__wctype "���  ___imp__pwctype "���  short int ܈  tm $"Q
��  
tm_sec "R	h   
tm_min "S	`      h  
tm_hour "T	h  
tm_mday "U	h  
tm_mon "V	h  
tm_year "W	h  
tm_wday "X	h  
tm_yday "Y	h  
tm_isdst "Z	h    �  mbstate_t "�h  ��  `btowc "�-  ҉  h   `fgetwc "-  �  �   ��  `fgetws "�  �  �  h  �   `fputwc "-  5�  �  �   `fputws "h  T�  T�  �   �  `fwide "�h  x�  �  h   afwprintf "Ih  ��  �  T�  b afwscanf "%h  ��  �  T�  b `getwc "-  Ԋ  �   cgetwchar "-  `mbrlen "��   
�  
�  �   �   �   
�  ��  `mbrtowc "��   E�  �  
�  �   �   `mbsinit "�h  `�  `�   ��  `mbsrtowcs "��   ��  �  ��  �   �   
�  `putwc "	-  ��  �  �   `putwchar "
-  ҋ  �   dp  #>h  �  �  T�  b dp  #"h  �  �  �   T�  b aswscanf "h  0�  T�  T�  b `ungetwc "-  P�  -  �   avfwprintf "_h  w�  �  T�  �    avfwscanf "?h  ��  �  T�  �    d
   #3h  ��  �  T�  �    d
   #h  �  �  �   T�  �    avswscanf "1h  �  T�  T�  �    avwprinta      f "fh  )�  T�  �    avwscanf "8h  I�  T�  �    `wcrtomb "��   n�  �  �  �   ewcscat $��  ��  �  T�   ewcscmp $�h  ��  T�  T�   ewcscoll $�h  ɍ  T�  T�   ewcscpy $��  �  �  T�   ewcscspn $��   �  T�  T�   `wcsftime "e�   1�  �  �   T�  1�   ��  ewcslen $��   P�  T�   ewcsncat $��  t�  �  T�  �    ewcsncmp $�h  ��  T�  T�  �    ewcsncpy $��  ��  �  T�  �    `wcsrtombs "��   �  �  �  �   �   T�  ewcsspn $��   �  T�  T�   awcstod "�+�  +�  T�  5�   double �  awcstof "�Z�  Z�  T�  5�   float ewcstok $��  ��  �  T�   `wcstol "�t  ��  T�  5�  h   `wcstoul "��  ʏ  T�  5�  h   ewcsxfrm $��   �  �  T�  �    `wctob "�h  �  -   `wmemcmp "�h  ,�  T�  T�  �    `wmemcpy "��  Q�  �  T�  �    `wmemmove "��  w�  �  T�  �    `wmemset "��  ��  �  �  �    awprintf "Th  ��  T�  b awscanf "h  Ӑ  T�  b ewcschr $�"�  �  T�  �   ewcspbrk $�"�  �  T�b        T�   ewcsrchr $�"�  /�  T�  �   ewcsstr $�"�  M�  T�  T�   `wmemchr "�"�  r�  T�  �  �    `wcstold "���  ��  T�  5�   long double `wcstoll "�'�   Ƒ  T�  5�  h   `wcstoull "�0�   �  T�  5�  h   �P  fjQ  �U  g�U  hdecltype(nullptr) ijQ  gjQ  bool %�  bV  2W   X  signed char �X  j Y  6__gnu_debug 8{�  P:>Y   g�Y  g�Y  �Y  �Y  g\  gf]  gs]  s]  f]  g�_  int8_t %#D�  uint8_t %$�  int16_t %%܈  uint16_t %&<  int32_t %'h  uint32_t %(�  int64_t %)&�   uint64_t %*0�   int_least8_t %-D�  uint_least8_t %.�  int_least16_t %/܈  uint_least16_t %0<  int_least32_t %1h  uint_least32_t %2�  int_least64_t %3&�   uint_least64_t %40�   int_fast8_t %:D�  uint_fast8_t %;�  int_fast16_t %<܈  uint_fast16_t %=<  int_fast32_t %>h  uint_fast32_t %?�  int_fast64_t %@&�   uint_fast64_t %A0�   intmax_t %D&�   uintmax_t %E0�   char16_t char32_t fpos_t &h%�   Д  esetlocale P�  �  h  c      
�   klocaleconv Q!�  �  #�  l ___newclmap 'P�  ___newcumap 'Q�  ___ptlocinfo 'R�  ___ptmbcinfo 'S�  ___globallocalestatus 'Th  ___locale_changed 'Uh  ___initiallocinfo 'V(�  ___initiallocalestructinfo 'W  ___imp___mb_cur_max '��  �  m
�  n�  h   ___security_cookie (}  n:�  �   /�  o_pthread_key_dest )#[�  :�  _Atomic_word * h  |�  p�n  g�q  �q  g�   g�   �a  gib  _div_t +;Ӗ  quot +<	h   rem +=	h   div_t +>��  _ldiv_t +@�  quot +A
t   rem +B
t   ldiv_t +C�  �  -�  �     __sys_errlist +�&�  __sys_nerr +�$h  o__imp___argc +�  o__imp___argv +��  ��  �  o__imp___wargv +!��  5�  o__imp__environ +'��  o__imp__wenviron +,��  o__imp__pgmptr +2��  o__imp__wpgmptr +75�  o__imp__osplatform +<$�  �  o__imp__osver +A$�  o__imp__winver +F$�  o__imp__winmajor +K$�  o__imp__winminor +P$�  q+�7lldiv_t ��  
quot +�0�    
rem +�6�    lldiv_t +�=��  __amblksiz ,5�  `atexit +�h  ��  ��   `d      atof +�+�  �  
�   `atoi +�h  '�  
�   `atol +�t  ?�  
�   `bsearch +��  n�  v�  v�  �   �   n�   t�  rh  ��  v�  v�   `div +�Ӗ  ��  h  h   `getenv +��  ��  
�   `ldiv +��  ۙ  t  t   `mblen +�h  ��  
�  �    `mbstowcs +��   �  �  
�  �    `mbtowc +�h  C�  �  
�  �    sqsort +�g�  �  �   �   n�   crand +�h  ssrand +���  �   astrtod +� +�  ��  
�  ��   `strtol +�t  ͚  
�  ��  h   `strtoul +��  �  
�  ��  h   esystem (Uh  �  
�   `wcstombs +��   1�  �  T�  �    `wctomb +�h  P�  �  �   `lldiv +�%��  n�  �   �    `atoll +�(�   ��  
�   `strtoll +�(�   ��  
�  ��  h   `strtoull +�1�   қ  
�  ��  h   astrtof +�Z�  �  
�  ��   `strtold +�'��  �  
�  ��   sclearerr &B)�  �   `fclose &Ch  C�  �   `feof &Jh  [�  �   `ferror &Kh  u�  �   `fflush &Lh  ��  �   `fgetc &Mh  ��  �   `fgetpos &Oh  Ȝ  �  Ȝ   Д  `fgets &Q�  �  �  h  �  e       `fopen &X�  �  
�  
�   afprintf &Nh  0�  �  
�  b `fread &]�   X�  �  �   �   �   `freopen &^�  }�  
�  
�  �   afscanf &!h  ��  �  
�  b `fseek &ah  ��  �  t  h   `fsetpos &_h  ��  �  ��   ߔ  `ftell &bt  ��  �   `getc &�h  �  �   cgetchar &�h  `gets &��  @�  �   sperror &�V�  
�   aprintf &Yh  q�  
�  b eremove -�h  ��  
�   erename -�h  ��  
�  
�   srewind &���  �   ascanf &h  ؞  
�  b ssetbuf &��  �  �   `setvbuf &�h  �  �  �  h  �    asprintf &dh  >�  �  
�  b asscanf &h  ^�  
�  
�  b ctmpfile &��  `tmpnam &��  ��  �   `ungetc &�h  ��  h  �   avfprintf &oh  Ο  �  
�  �    avprintf &vh  �  
�  �    avsprintf &}h  �  �  
�  �    asnprintf &�h  ;�  �  �   
�  b avfscanf &@h  `�  �  
�  �    avscanf &9h  �  
�  �    avsnprintf &�h  ��  �  �   
�  �    avsscanf &2h  Р  
�  
�  �    g7e  gDe  g�a  gfu  f      gru  a  i�a  �   
�  �      �N  g�  gM  gZ  g�N  i  g  g  �h  �i  wctrans_t .��  `iswctype "#h  �  -  W   etowctrans .�-  ��  -  L�   ewctrans .�L�  ��  
�   ewctype .�W  ӡ  
�   t�l  	0�L     _PHNDLR /?�  _XCPT_ACTION /A
>�  XcptNum /B�   SigNum /C	h  XcptAction /D�   �  I�  l __XcptActTab /G>�  __XcptActTabCount /Hh  __XcptActTabSize /Ih  __First_FPE_Indx /Jh  __Num_FPE /Kh  DWORD 0��  _GUID 1�  Data1 1�   Data2 1<  Data3 1<  Data4 1�   �  !�  �    GUID 1Ţ  !�  IID 1S!�  3�  CLSID 1[!�  D�  FMTID 1b!�  W�  oGUID_MAX_POWER_SAVINGS 2�.�  oGUID_MIN_POWER_SAVINGS 2�.�  oGUID_TYPICAL_POWER_SAVINGS 2�.�  oNO_SUBGROUP_GUID 2�.�  oALL_POWERSCHEMES_GUID 2�.�  oGUID_POWERSCHEME_PERSONALITY 2�.�  oGUID_ACTIVE_POWERSCHEME 2�.�  oGUID_IDLE_RESILIENCY_SUBGROUP 2�.�  oGUID_IDLE_RESILIENCY_PERIOD 2�.�  oGUID_DISK_COALESCING_POWERDOWN_TIMEOUT 2�.�  oGUID_EXECUTION_REQUIRg      ED_REQUEST_TIMEOUT 2�.�  oGUID_VIDEO_SUBGROUP 2�.�  oGUID_VIDEO_POWERDOWN_TIMEOUT 2�.�  oGUID_VIDEO_ANNOYANCE_TIMEOUT 2�.�  oGUID_VIDEO_ADAPTIVE_PERCENT_INCREASE 2�.�  oGUID_VIDEO_DIM_TIMEOUT 2�.�  oGUID_VIDEO_ADAPTIVE_POWERDOWN 2�.�  oGUID_MONITOR_POWER_ON 2�.�  oGUID_DEVICE_POWER_POLICY_VIDEO_BRIGHTNESS 2�.�  oGUID_DEVICE_POWER_POLICY_VIDEO_DIM_BRIGHTNESS 2�.�  oGUID_VIDEO_CURRENT_MONITOR_BRIGHTNESS 2�.�  oGUID_VIDEO_ADAPTIVE_DISPLAY_BRIGHTNESS 2�.�  oGUID_CONSOLE_DISPLAY_STATE 2�.�  oGUID_ALLOW_DISPLAY_REQUIRED 2�.�  oGUID_VIDEO_CONSOLE_LOCK_TIMEOUT 2�.�  oGUID_ADAPTIVE_POWER_BEHAVIOR_SUBGROUP 2�.�  oGUID_NON_ADAPTIVE_INPUT_TIMEOUT 2�.�  oGUID_DISK_SUBGROUP 2�.�  oGUID_DISK_POWERDOWN_TIMEOUT 2�.�  oGUID_DISK_IDLE_TIMEOUT 2�.�  oGUID_DISK_BURST_IGNORE_THRESHOLD 2�.�  oGUID_DISK_ADAPTIVE_POWERDOWN 2�.�  oGUID_SLEEP_SUBGROUP 2�.�  oGUID_SLEEP_IDLE_THRESHOLD 2�.�  oGUID_STANDBY_TIMEOUT 2�.�  oGUID_UNATTEND_SLEEP_TIMEOUT 2�.�  oGUID_HIBERNATE_TIMEOUT 2h      �.�  oGUID_HIBERNATE_FASTS4_POLICY 2�.�  oGUID_CRITICAL_POWER_TRANSITION 2�.�  oGUID_SYSTEM_AWAYMODE 2�.�  oGUID_ALLOW_AWAYMODE 2�.�  oGUID_ALLOW_STANDBY_STATES 2�.�  oGUID_ALLOW_RTC_WAKE 2�.�  oGUID_ALLOW_SYSTEM_REQUIRED 2�.�  oGUID_SYSTEM_BUTTON_SUBGROUP 2�.�  oGUID_POWERBUTTON_ACTION 2�.�  oGUID_SLEEPBUTTON_ACTION 2�.�  oGUID_USERINTERFACEBUTTON_ACTION 2�.�  oGUID_LIDCLOSE_ACTION 2�.�  oGUID_LIDOPEN_POWERSTATE 2�.�  oGUID_BATTERY_SUBGROUP 2�.�  oGUID_BATTERY_DISCHARGE_ACTION_0 2�.�  oGUID_BATTERY_DISCHARGE_LEVEL_0 2�.�  oGUID_BATTERY_DISCHARGE_FLAGS_0 2�.�  oGUID_BATTERY_DISCHARGE_ACTION_1 2�.�  oGUID_BATTERY_DISCHARGE_LEVEL_1 2�.�  oGUID_BATTERY_DISCHARGE_FLAGS_1 2�.�  oGUID_BATTERY_DISCHARGE_ACTION_2 2�.�  oGUID_BATTERY_DISCHARGE_LEVEL_2 2�.�  oGUID_BATTERY_DISCHARGE_FLAGS_2 2�.�  oGUID_BATTERY_DISCHARGE_ACTION_3 2�.�  oGUID_BATTERY_DISCHARGE_LEVEL_3 2�.�  oGUID_BATTERY_DISCHARGE_FLAGS_3 2�.�  oGUID_PROCESSOR_SETTINGS_SUBGROUP 2�.�  oGUID_PRi      OCESSOR_THROTTLE_POLICY 2�.�  oGUID_PROCESSOR_THROTTLE_MAXIMUM 2�.�  oGUID_PROCESSOR_THROTTLE_MINIMUM 2�.�  oGUID_PROCESSOR_ALLOW_THROTTLING 2�.�  oGUID_PROCESSOR_IDLESTATE_POLICY 2�.�  oGUID_PROCESSOR_PERFSTATE_POLICY 2�.�  oGUID_PROCESSOR_PERF_INCREASE_THRESHOLD 2�.�  oGUID_PROCESSOR_PERF_DECREASE_THRESHOLD 2�.�  oGUID_PROCESSOR_PERF_INCREASE_POLICY 2�.�  oGUID_PROCESSOR_PERF_DECREASE_POLICY 2�.�  oGUID_PROCESSOR_PERF_INCREASE_TIME 2�.�  oGUID_PROCESSOR_PERF_DECREASE_TIME 2�.�  oGUID_PROCESSOR_PERF_TIME_CHECK 2�.�  oGUID_PROCESSOR_PERF_BOOST_POLICY 2�.�  oGUID_PROCESSOR_PERF_BOOST_MODE 2�.�  oGUID_PROCESSOR_IDLE_ALLOW_SCALING 2�.�  oGUID_PROCESSOR_IDLE_DISABLE 2�.�  oGUID_PROCESSOR_IDLE_STATE_MAXIMUM 2�.�  oGUID_PROCESSOR_IDLE_TIME_CHECK 2�.�  oGUID_PROCESSOR_IDLE_DEMOTE_THRESHOLD 2�.�  oGUID_PROCESSOR_IDLE_PROMOTE_THRESHOLD 2�.�  oGUID_PROCESSOR_CORE_PARKING_INCREASE_THRESHOLD 2�.�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_THRESHOLD 2�.�  oGUID_PROCESSOR_Cj      ORE_PARKING_INCREASE_POLICY 2 .�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_POLICY 2.�  oGUID_PROCESSOR_CORE_PARKING_MAX_CORES 2.�  oGUID_PROCESSOR_CORE_PARKING_MIN_CORES 2.�  oGUID_PROCESSOR_CORE_PARKING_INCREASE_TIME 2.�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_TIME 2.�  oGUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_DECREASE_FACTOR 2.�  oGUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_THRESHOLD 2.�  oGUID_PROCESSOR_CORE_PARKING_AFFINITY_WEIGHTING 2.�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_DECREASE_FACTOR 2	.�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_THRESHOLD 2
.�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_WEIGHTING 2.�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_THRESHOLD 2.�  oGUID_PROCESSOR_PARKING_CORE_OVERRIDE 2.�  oGUID_PROCESSOR_PARKING_PERF_STATE 2.�  oGUID_PROCESSOR_PARKING_CONCURRENCY_THRESHOLD 2.�  oGUID_PROCESSOR_PARKING_HEADROOM_THRESHOLD 2.�  oGUID_PROCESSOR_PERF_HISTORY 2.�  oGUID_PROCESSOR_PERF_LATENCY_HINk      T 2.�  oGUID_PROCESSOR_DISTRIBUTE_UTILITY 2.�  oGUID_SYSTEM_COOLING_POLICY 2.�  oGUID_LOCK_CONSOLE_ON_WAKE 2.�  oGUID_DEVICE_IDLE_POLICY 2.�  oGUID_ACDC_POWER_SOURCE 2.�  oGUID_LIDSWITCH_STATE_CHANGE 2.�  oGUID_BATTERY_PERCENTAGE_REMAINING 2.�  oGUID_GLOBAL_USER_PRESENCE 2.�  oGUID_SESSION_DISPLAY_STATUS 2.�  oGUID_SESSION_USER_PRESENCE 2.�  oGUID_IDLE_BACKGROUND_TASK 2.�  oGUID_BACKGROUND_TASK_NOTIFICATION 2.�  oGUID_APPLAUNCH_BUTTON 2.�  oGUID_PCIEXPRESS_SETTINGS_SUBGROUP 2 .�  oGUID_PCIEXPRESS_ASPM_POLICY 2!.�  oGUID_ENABLE_SWITCH_FORCED_SHUTDOWN 2".�  oPPM_PERFSTATE_CHANGE_GUID 2 .�  oPPM_PERFSTATE_DOMAIN_CHANGE_GUID 2!.�  oPPM_IDLESTATE_CHANGE_GUID 2".�  oPPM_PERFSTATES_DATA_GUID 2#.�  oPPM_IDLESTATES_DATA_GUID 2$.�  oPPM_IDLE_ACCOUNTING_GUID 2%.�  oPPM_IDLE_ACCOUNTING_EX_GUID 2&.�  oPPM_THERMALCONSTRAINT_GUID 2'.�  oPPM_PERFMON_PERFSTATE_GUID 2(.�  oPPM_THERMAL_POLICY_CHANGE_GUID 2).�  RPC_IF_HANDLE 3B�  24'ݘ  243Ӗ  244l      �  `abs +h  Ҹ  h   246��  246m  246,m  246Lm  246lm  246�m  247��  248�  249'�  24:?�  24<*r  24<��  24<�m  24>��  24@��  24Cۙ  24D��  24E�  24GC�  24Hg�  24Ju�  24K��  24L��  24M͚  24N�  24P�  24Q1�  _IWinTypesBase_v0_1_c_ifspec 5)��  _IWinTypesBase_v0_1_s_ifspec 5*��  _IID_IUnknown 6=?�  _IID_AsyncIUnknown 6�.�  oIID_IClassFactory 6m.�  oIID_IMarshal 7n.�  oIID_INoMarshal 7U.�  oIID_IAgileObject 7�.�  oIID_IAgileReference 7�.�  oIID_IMarshal2 7-.�  oIID_IMalloc 7�.�  oIID_IStdMarshalInfo 7i.�  oIID_IExternalConnection 7�.�  oIID_IMultiQI 7G.�  oIID_AsyncIMultiQI 7�.�  oIID_IInternalUnknown 7.�  oIID_IEnumUnknown 7h.�  oIID_IEnumString 7.�  oIID_ISequentialStream 7�.�  oIID_IStream 7M.�  oIID_IRpcChannelBuffer 7�	.�  oIID_IRpcChannelBuffer2 7;
.�  oIID_IAsyncRpcChannelBuffer 7�
.�  oIID_IRpcChannelBuffer3 7.�  oIID_IRpcSyntaxNegotiate 7�.�  oIID_IRpcProxyBuffer 7�.�  oIID_IRpcStubBuffer 7V.�  oIID_IPSFactoryBufm      fer 7.�  oIID_IChannelHook 7�.�  oIID_IClientSecurity 7�.�  oIID_IServerSecurity 7m.�  oIID_IRpcOptions 7.�  oIID_IGlobalOptions 7�.�  oIID_ISurrogate 7!.�  oIID_IGlobalInterfaceTable 7�.�  oIID_ISynchronize 7.�  oIID_ISynchronizeHandle 7�.�  oIID_ISynchronizeEvent 7�.�  oIID_ISynchronizeContainer 7A.�  oIID_ISynchronizeMutex 7�.�  oIID_ICancelMethodCalls 7.�  oIID_IAsyncManager 7�.�  oIID_ICallFactory 7.�  oIID_IRpcHelper 7f.�  oIID_IReleaseMarshalBuffers 7�.�  oIID_IWaitMultiple 7,.�  oIID_IAddrTrackingControl 7�.�  oIID_IAddrExclusionControl 7�.�  oIID_IPipeByte 7h.�  oIID_IPipeLong 7�.�  oIID_IPipeDouble 7J.�  oIID_IComThreadingInfo 7$.�  oIID_IProcessInitControl 7�.�  oIID_IFastRundown 7.�  oIID_IMarshalingStream 7J.�  oIID_ICallbackWithNoReentrancyToApplicationSTA 7	.�  _GUID_NULL 8?�  _CATID_MARSHALER 8?�  _IID_IRpcChannel 8?�  _IID_IRpcStub 8?�  _IID_IStubManager 8?�  _IID_IRpcProxy 8?�  _IID_IProxyManager 8?�  _IID_n      IPSFactory 8?�  _IID_IInternalMoniker 8?�  _IID_IDfReserved1 8?�  _IID_IDfReserved2 8?�  _IID_IDfReserved3 8?�  _CLSID_StdMarshal 8R�  _CLSID_AggStdMarshal 8R�  _CLSID_StdAsyncActManager 8R�  _IID_IStub 8?�  _IID_IProxy 8?�  _IID_IEnumGeneric 8?�  _IID_IEnumHolder 8?�  _IID_IEnumCallback 8 ?�  _IID_IOleManager 8!?�  _IID_IOlePresObj 8"?�  _IID_IDebug 8#?�  _IID_IDebugStream 8$?�  _CLSID_PSGenObject 8%R�  _CLSID_PSClientSite 8&R�  _CLSID_PSClassObject 8'R�  _CLSID_PSInPlaceActive 8(R�  _CLSID_PSInPlaceFrame 8)R�  _CLSID_PSDragDrop 8*R�  _CLSID_PSBindCtx 8+R�  _CLSID_PSEnumerators 8,R�  _CLSID_StaticMetafile 8-R�  _CLSID_StaticDib 8.R�  _CID_CDfsVolume 8/R�  _CLSID_DCOMAccessControl 80R�  _CLSID_GlobalOptions 81R�  _CLSID_StdGlobalInterfaceTable 82R�  _CLSID_ComBinding 83R�  _CLSID_StdEvent 84R�  _CLSID_ManualResetEvent 85R�  _CLSID_SynchronizeContainer 86R�  _CLSID_AddrControl 87R�  _CLSID_CCDFormKrnl 88R�  _CLSID_CCDPropertyPage 89R�  _CLSID_CCDFormDiao      log 8:R�  _CLSID_CCDCommandButton 8;R�  _CLSID_CCDComboBox 8<R�  _CLSID_CCDTextBox 8=R�  _CLSID_CCDCheckBox 8>R�  _CLSID_CCDLabel 8?R�  _CLSID_CCDOptionButton 8@R�  _CLSID_CCDListBox 8AR�  _CLSID_CCDScrollBar 8BR�  _CLSID_CCDGroupBox 8CR�  _CLSID_CCDGeneralPropertyPage 8DR�  _CLSID_CCDGenericPropertyPage 8ER�  _CLSID_CCDFontPropertyPage 8FR�  _CLSID_CCDColorPropertyPage 8GR�  _CLSID_CCDLabelPropertyPage 8HR�  _CLSID_CCDCheckBoxPropertyPage 8IR�  _CLSID_CCDTextBoxPropertyPage 8JR�  _CLSID_CCDOptionButtonPropertyPage 8KR�  _CLSID_CCDListBoxPropertyPage 8LR�  _CLSID_CCDCommandButtonPropertyPage 8MR�  _CLSID_CCDComboBoxPropertyPage 8NR�  _CLSID_CCDScrollBarPropertyPage 8OR�  _CLSID_CCDGroupBoxPropertyPage 8PR�  _CLSID_CCDXObjectPropertyPage 8QR�  _CLSID_CStdPropertyFrame 8RR�  _CLSID_CFormPropertyPage 8SR�  _CLSID_CGridPropertyPage 8TR�  _CLSID_CWSJArticlePage 8UR�  _CLSID_CSystemPage 8VR�  _CLSID_IdentityUnmarshal 8WR�  _CLSID_InProcFreeMarshaler 8XR�  _CLSID_Picture_Metafip      le 8YR�  _CLSID_Picture_EnhMetafile 8ZR�  _CLSID_Picture_Dib 8[R�  _GUID_TRISTATE 8\.�  _IWinTypes_v0_1_c_ifspec 9(��  _IWinTypes_v0_1_s_ifspec 9)��  oIID_IMallocSpy :�.�  oIID_IBindCtx ::.�  oIID_IEnumMoniker :J .�  oIID_IRunnableObject :� .�  oIID_IRunningObjectTable :�!.�  oIID_IPersist :i".�  oIID_IPersistStream :�".�  oIID_IMoniker :j#.�  oIID_IROTData :X%.�  oIID_IEnumSTATSTG :�%.�  oIID_IStorage :X&.�  oIID_IPersistFile :A(.�  oIID_IPersistStorage :�(.�  oIID_ILockBytes :�).�  oIID_IEnumFORMATETC :�*.�  oIID_IEnumSTATDATA :l+.�  oIID_IRootStorage :,.�  oIID_IAdviseSink :�,.�  oIID_AsyncIAdviseSink :s-.�  oIID_IAdviseSink2 :�..�  oIID_AsyncIAdviseSink2 :./.�  oIID_IDataObject :�/.�  oIID_IDataAdviseHolder :1.�  oIID_IMessageFilter :�1.�  oFMTID_SummaryInformation :]2e�  oFMTID_DocSummaryInformation :_2e�  oFMTID_UserDefinedProperties :a2e�  oFMTID_DiscardableInformation :c2e�  oFMTID_ImageSummaryInformation :e2e�  oFMTID_AudioSummaryInformation :g2e�  oFMTq      ID_VideoSummaryInformation :i2e�  oFMTID_MediaFileSummaryInformation :k2e�  oIID_IClassActivator :s2.�  oIID_IFillLockBytes :�2.�  oIID_IProgressNotify :�3.�  oIID_ILayoutStorage :�3.�  oIID_IBlockingLock :�4.�  oIID_ITimeAndNoticeControl :�4.�  oIID_IOplockStorage :N5.�  oIID_IDirectWriterLock :�5.�  oIID_IUrlMon :M6.�  oIID_IForegroundTransfer :�6.�  oIID_IThumbnailExtractor :7.�  oIID_IDummyHICONIncluder :�7.�  oIID_IProcessLock :�7.�  oIID_ISurrogateService :H8.�  oIID_IInitializeSpy :�8.�  oIID_IApartmentShutdown :�9.�  _IID_IOleAdviseHolder ;�.�  oIID_IOleCache ;b.�  oIID_IOleCache2 ;).�  oIID_IOleCacheControl ;�.�  oIID_IParseDisplayName ;<.�  oIID_IOleContainer ;�.�  oIID_IOleClientSite ;.�  oIID_IOleObject ;�.�  oIOLETypes_v0_0_c_ifspec ;���  oIOLETypes_v0_0_s_ifspec ;���  oIID_IOleWindow ;$.�  oIID_IOleLink ;�.�  oIID_IOleItemContainer ;�.�  oIID_IOleInPlaceUIWindow ;v	.�  oIID_IOleInPlaceActiveObject ;
.�  oIID_IOleInPlaceFrame ;�
.�  oIID_IOr      leInPlaceObject ;�.�  oIID_IOleInPlaceSite ;�.�  oIID_IContinue ;�.�  oIID_IViewObject ;�.�  oIID_IViewObject2 ;*.�  oIID_IDropSource ;�.�  oIID_IDropTarget ;[.�  oIID_IDropSourceNotify ;�.�  oIID_IEnumOLEVERB ;v.�  _IID_IServiceProvider <9?�  _IOleAutomationTypes_v1_0_c_ifspec =���  _IOleAutomationTypes_v1_0_s_ifspec =���  oIID_ICreateTypeInfo =;.�  oIID_ICreateTypeInfo2 =b.�  oIID_ICreateTypeLib =�.�  oIID_ICreateTypeLib2 =�.�  oIID_IDispatch =�	.�  oIID_IEnumVARIANT =�
.�  oIID_ITypeComp =5.�  oIID_ITypeInfo =�.�  oIID_ITypeInfo2 =P.�  oIID_ITypeLib =�.�  oIID_ITypeLib2 ==.�  oIID_ITypeChangeEvents =a.�  oIID_IErrorInfo =�.�  oIID_ICreateErrorInfo =}.�  oIID_ISupportErrorInfo = .�  oIID_ITypeFactory =u.�  oIID_ITypeMarshal =�.�  oIID_IRecordInfo =�.�  oIID_IErrorLog = .�  oIID_IPropertyBag =z.�  ___MIDL_itf_msxml_0000_v0_0_c_ifspec >���  ___MIDL_itf_msxml_0000_v0_0_s_ifspec >���  _LIBID_MSXML >�?�  oIID_IXMLDOMImplementation > ?�  oIIDs      _IXMLDOMNode >'?�  oIID_IXMLDOMDocumentFragment >�?�  oIID_IXMLDOMDocument >f?�  oIID_IXMLDOMNodeList >u?�  oIID_IXMLDOMNamedNodeMap >�?�  oIID_IXMLDOMCharacterData >?�  oIID_IXMLDOMAttribute >�?�  oIID_IXMLDOMElement >?�  oIID_IXMLDOMText >�?�  oIID_IXMLDOMComment >%?�  oIID_IXMLDOMProcessingInstruction >�?�  oIID_IXMLDOMCDATASection >?�  oIID_IXMLDOMDocumentType >�?�  oIID_IXMLDOMNotation >?�  oIID_IXMLDOMEntity >?�  oIID_IXMLDOMEntityReference >�?�  oIID_IXMLDOMParseError >a	?�  oIID_IXTLRuntime >�	?�  oDIID_XMLDOMDocumentEvents >=
?�  oCLSID_DOMDocument >\
R�  oCLSID_DOMFreeThreadedDocument >`
R�  oIID_IXMLHttpRequest >g
?�  oCLSID_XMLHTTPRequest >�
R�  oIID_IXMLDSOControl >�
?�  oCLSID_XMLDSOControl >R�  oIID_IXMLElementCollection >?�  oIID_IXMLDocument >J?�  oIID_IXMLDocument2 >�?�  oIID_IXMLElement >$?�  oIID_IXMLElement2 >�?�  oIID_IXMLAttribute >�?�  oIID_IXMLError >?�  oCLSID_XMLDocument >.R�  oCLSID_SBS_StdURLMoniker ?~?�  t      oCLSID_SBS_HttpProtocol ??�  oCLSID_SBS_FtpProtocol ?�?�  oCLSID_SBS_GopherProtocol ?�?�  oCLSID_SBS_HttpSProtocol ?�?�  oCLSID_SBS_FileProtocol ?�?�  oCLSID_SBS_MkProtocol ?�?�  oCLSID_SBS_UrlMkBindCtx ?�?�  oCLSID_SBS_SoftDistExt ?�?�  oCLSID_SBS_CdlProtocol ?�?�  oCLSID_SBS_ClassInstallFilter ?�?�  oCLSID_SBS_InternetSecurityManager ?�?�  oCLSID_SBS_InternetZoneManager ?�?�  oIID_IAsyncMoniker ?�?�  oCLSID_StdURLMoniker ?�?�  oCLSID_HttpProtocol ?�?�  oCLSID_FtpProtocol ?�?�  oCLSID_GopherProtocol ?�?�  oCLSID_HttpSProtocol ?�?�  oCLSID_FileProtocol ?�?�  oCLSID_MkProtocol ?�?�  oCLSID_StdURLProtocol ?�?�  oCLSID_UrlMkBindCtx ?�?�  oCLSID_CdlProtocol ?�?�  oCLSID_ClassInstallFilter ?�?�  oIID_IAsyncBindCtx ?�?�  oIID_IPersistMoniker ?P.�  oIID_IMonikerProp ?!.�  oIID_IBindProtocol ?.�  oIID_IBinding ?�.�  oIID_IBindStatusCallback ?u.�  oIID_IBindStatusCallbackEx ?�.�  oIID_IAuthenticate ?d.�  oIID_IAuthenticateEx ?�.�  oIID_IHttpNeu      gotiate ?A.�  oIID_IHttpNegotiate2 ?�.�  oIID_IHttpNegotiate3 ?;	.�  oIID_IWinInetFileStream ?�	.�  oIID_IWindowForBindingUI ?0
.�  oIID_ICodeInstall ?�
.�  oIID_IWinInetInfo ?�.�  oIID_IHttpSecurity ?.�  oIID_IWinInetHttpInfo ?y.�  oIID_IWinInetHttpTimeouts ?�.�  oSID_BindHost ?5.�  oIID_IBindHost ??.�  oIID_IInternet ?M.�  oIID_IInternetBindInfo ?�.�  oIID_IInternetBindInfoEx ?&.�  oIID_IInternetProtocolRoot ?�.�  oIID_IInternetProtocol ?�.�  oIID_IInternetProtocolSink ?.�  oIID_IInternetProtocolSinkStackable ?�.�  oIID_IInternetSession ??.�  oIID_IInternetThreadSwitch ?H.�  oIID_IInternetPriority ?�.�  oIID_IInternetProtocolInfo ?N.�  oCLSID_InternetSecurityManager ?�?�  oCLSID_InternetZoneManager ?�?�  oIID_IInternetSecurityMgrSite ?�.�  oIID_IInternetSecurityManager ?i.�  oIID_IInternetHostSecurityManager ?!.�  oIID_IInternetZoneManager ?�".�  oCLSID_SoftDistExt ?�&?�  oIID_ISoftDistExt ?�&.�  oIID_ICatalogFileInfo ?x'.�  oIID_IDataFilter v      ?�'.�  oIID_IEncodingFilterFactory ?�(.�  oGUID_CUSTOM_CONFIRMOBJECTSAFETY ?3).�  oIID_IWrappedProtocol ?A).�  oIID_IGetBindHandle ?�).�  oIID_IBindCallbackRedirect ?*.�  oIID_IPropertyStorage @�.�  oIID_IPropertySetStorage @.�  oIID_IEnumSTATPROPSTG @�.�  oIID_IEnumSTATPROPSETSTG @D.�  _IID_StdOle A?�  _GUID_DEVINTERFACE_DISK B.�  _GUID_DEVINTERFACE_CDROM B.�  _GUID_DEVINTERFACE_PARTITION B.�  _GUID_DEVINTERFACE_TAPE B.�  _GUID_DEVINTERFACE_WRITEONCEDISK B.�  _GUID_DEVINTERFACE_VOLUME B.�  _GUID_DEVINTERFACE_MEDIUMCHANGER B.�  _GUID_DEVINTERFACE_FLOPPY B.�  _GUID_DEVINTERFACE_CDCHANGER B.�  _GUID_DEVINTERFACE_STORAGEPORT B.�  _GUID_DEVINTERFACE_COMPORT B.�  _GUID_DEVINTERFACE_SERENUM_BUS_ENUMERATOR B.�  _SCARD_IO_REQUEST C���  dwProtocol C���   cbPciLength C���   SCARD_IO_REQUEST C�\�  ��  _g_rgSCardT0Pci D%.��  _g_rgSCardT1Pci D%=��  _g_rgSCardRawPci D%L��  _IID_IPrintDialogCallback E.�  _IID_IPrintDialogServices E.�  2F�N  2F2l  }}  gw      �  �  g}}  �u  g�  x}  g�u  u_ZNSt17integral_constantIbLb0EE5valueE �V   u_ZNSt17integral_constantIbLb1EE5valueE ^W  v_ZN9__gnu_cxx24__numeric_traits_integerIiE5__minE �q  ����xw_ZN9__gnu_cxx24__numeric_traits_integerIiE5__maxE �q  ���u_ZN9__gnu_cxx25__numeric_traits_floatingIfE16__max_exponent10E q�  &x_ZN9__gnu_cxx25__numeric_traits_floatingIdE16__max_exponent10E օ  4x_ZN9__gnu_cxx25__numeric_traits_floatingIeE16__max_exponent10E @�  Du_ZN9__gnu_cxx24__numeric_traits_integerImE8__digitsE ��   u_ZN9__gnu_cxx24__numeric_traits_integerIcE5__maxE ��  v_ZN9__gnu_cxx24__numeric_traits_integerIsE5__minE T�  ��~x_ZN9__gnu_cxx24__numeric_traits_integerIsE5__maxE `�  �v_ZN9__gnu_cxx24__numeric_traits_integerIxE5__minE ��  ���������y_ZN9__gnu_cxx24__numeric_traits_integerIxE5__maxE Ǉ  �������z_GLOBAL__sub_I_main �@            �{__static_initialization_and_destruction_0 �@     <       �(�  |__initialize_p h  � |__priority h  � z__tcf_0 �@            �}main h  P@     x      ?       � H�     GNU C++11 8.1.0 -mtune=core2 -march=nocona -g -std=c++11 F:\debug\ClionWork\EFS\OS\VHD\disk.cpp F:\debug\ClionWork\EFS\cmake-build-debug @     u         __builtin_va_list �   char �   size_t #,�   long long unsigned int long long int �   intptr_t >#�   uintptr_t K,�   wint_t j@  short unsigned int @  wctype_t k@  int l  long int pthreadlocinfo �(�  �  threadlocaleinfostruct `��  	 �
  
locale ��   
wlocale ��  �  �
�  
wrefcount �
�   �  �l   
lc_codepage ��  
lc_collate_cp ��  
lc_handle ��  
lc_id ��  $
lc_category ��  Hlc_clike �l  mb_cur_max �l  lconv_intl_refcount ��  lconv_num_refcount ��  lconv_mon_refcount ��   lconv ��  (ctype1_refcount ��  0ctype1 ��  8pctype ��  @pclmap ��  Hpcumap ��  Plc_time_curr ��  X pthreadmbcinfo �%�  �  threadmbcinfostruct localeinfo_struct �  
ly      ocinfo ��   
mbcinfo ��   _locale_tstruct ��  tagLC_ID �x  
wLanguage �@   
wCountry �@  
wCodePage �@   LC_ID �)  �   �  �  wchar_t �  l  unsigned int �  �  �    long unsigned int �  x  �  �    �    �    lconv X-
�  decimal_point .�   thousands_sep /�  grouping 0�  int_curr_symbol 1�  currency_symbol 2�   mon_decimal_point 3�  (mon_thousands_sep 4�  0mon_grouping 5�  8positive_sign 6�  @negative_sign 7�  Hint_frac_digits 8
�   Pfrac_digits 9
�   Qp_cs_precedes :
�   Rp_sep_by_space ;
�   Sn_cs_precedes <
�   Tn_sep_by_space =
�   Up_sign_posn >
�   Vn_sign_posn ?
�   W   @  V  �  unsigned char �  __lc_time_data �  std G un  __cxx11 
A�N  basic_string<char, std::char_traits<char>, std::allocator<char> >  M�N  7  �b  �a   7  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC4EPcRKS3_ �  �  �  b  ��  z       7  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC4EPcOS3_ C  S  �  b  ��   _M_p �
b    �  \0{u  ��  _M_local_buf �5��  _M_allocated_capacity ��     X2�u  �  npos e�  _M_dataplus �e   _M_string_length ��  o   _M_data �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc V	  a	  �  b    _M_length �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy �	  �	  �  �   !_M_data �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv b  
  #
  �   "J  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv b  ~
  �
  �   �  ]5�u  "J  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv �
  �
  �
  �    _M_capacity �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy P  [  �  �    _M_set_length �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy �  �  �  �   !_M_is_local �_ZNKSt{      7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv )�  )  /  �   !_M_create �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy b  �  �  �  �  �    _M_dispose �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv �  �  �    _M_destroy �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy Y  d  �  �    _M_construct_aux_2 �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc �  �  �  �  �    #_M_construct _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructEyc A  Q  �  �  �      W#c  Q  _Char_alloc_type P�u  $q  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv  �  �  �  �   $q  _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv &�  A  G  �   %_M_check +_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc �  �  �  �  �  �   #_M_check_length 5_ZNKSt7__c|      xx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc !  6  �  �  �  �   %_M_limit >_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy �  �  �  �  �  �   %_M_disjunct F_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc )�      �  �   &_S_copy O_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy y  �  �  �   &_S_move X_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy �  �  �  �   &_S_assign a_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_S_assignEPcyc G  �  �  �    '#  t_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ �  �  �  �   �  ^D�u  '#  x_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcS4_EESA_ r  �  r  r   )  `�}  '#  }_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsE}      PcS5_S5_ �  �  �  �   '#  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ U  �  �  �   (_S_compare �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy l  �  �  �   #_M_assign �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_assignERKS4_   %  �  ,�   #_M_mutate �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy �  �  �  �  �  �  �   #_M_erase �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy �    �  �  �   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4Ev Q  W  �   *�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS3_ �  �  �  ��   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_     �  ,�   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yRKS3_ c  x  �  ,�  �  ��   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yy � ~       �  �  ,�  �  �   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_yyRKS3_ 6  P  �  ,�  �  �  ��   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EPKcyRKS3_ �  �  �  �  �  ��   )�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EPKcRKS3_     �  �  ��   )�  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EycRKS3_ n  �  �  �  �   ��   )�  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EOS4_ �  �  �  2�   )�  ._ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ESt16initializer_listIcERKS3_ D  T  �  g  ��   )�  2_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4ERKS4_RKS3_ �  �  �  ,�  ��   )�  6_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC4EOS4_RKS3_     �  2�  ��   +~basic_string �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED4Ei s  ~  �  l   ,|  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEa      SERKS4_ 8�  �  �  �  ,�   ,|  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEPKc 8�  /  :  �  �   ,|  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc 8�  �  �  �  �    ,|  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ 8�  �  �  �  2�   ,|  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE 8�  Y  d  �  g   -begin '_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv �  �  �  �   -begin /_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv r      �   -end 7_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv �  o  u  �   -end ?_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv r  �  �  �   .reverse_iterator b0�h  -rbegin H_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv �  @  F  �   .const_reverse_iterator a5Ri  -rbegin Q_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv F �       �  �  �   -rend Z_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv �        �   -rend c_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv F  t   z   �   -cbegin l_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv r  �   �   �   -cend t_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv r  .!  4!  �   -crbegin }_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv F  �!  �!  �   -crend �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv F  �!  �!  �   -size �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv �  G"  M"  �   ,h  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv �  �"  �"  �   ,�  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8max_sizeEv �  #  #  �   +resize �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc \#  l#  �  �  �    +resize �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE�      6resizeEy �#  �#  �  �   +shrink_to_fit �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv .$  4$  �   -capacity �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv �  �$  �$  �   +reserve �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy �$  �$  �  �   +clear �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv J%  P%  �   -empty �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv )�  �%  �%  �   d  [7�u  ,�  _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy �%  &  &  �  �   O  Z2�u  ,�  _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy &  s&  ~&  �  �   -at )_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy �%  �&  �&  �  �   -at >_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy &  *'  5'  �  �   -front N_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv &  �'  �'  �   -front Y_ZNKSt7__�      cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv �%  �'  �'  �   -back d_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv &  B(  H(  �   -back o_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv �%  �(  �(  �   ,  }_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ 8�  �(  )  �  ,�   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc 8�  T)  _)  �  �   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc 8�  �)  �)  �  �    ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE 8�   *  +*  �  g   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ 8�  �*  �*  �  ,�   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy 8�  �*  �*  �  ,�  �  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy 8�  W+  g+  �  �  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsI�      cESaIcEE6appendEPKc 8�  �+  �+  �  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc 8�  ,  /,  �  �  �    ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendESt16initializer_listIcE 8�  �,  �,  �  g   +push_back 2_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9push_backEc �,  
-  �  �    ,  A_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ 8�  c-  n-  �  ,�   ,  Q_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ 8�  �-  �-  �  2�   ,  h_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy 8�  ,.  A.  �  ,�  �  �   ,  x_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKcy 8�  �.  �.  �  �  �   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc 8�   /  /  �  �   ,  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc 8�  a/  q/  �  �  �    ,  �_ZNSt7__cxx1112basic_string�      IcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE 8�  �/  �/  �  g   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc �  d0  y0  �  r  �  �    )�  8_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE 1  1  �  �  g   ,�  L_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ 8�  p1  �1  �  �  ,�   ,�  c_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_yy 8�  �1  �1  �  �  ,�  �  �   ,�  z_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy 8�  O2  d2  �  �  �  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKc 8�  �2  �2  �  �  �   ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc 8�  #3  83  �  �  �  �    ,�  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__�      normal_iteratorIPKcS4_EEc �  �3  �3  �  �3  �    __const_iterator lr  -erase �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy 8�  44  D4  �  �  �   -erase _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE �  �4  �4  �  �3   -erase _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ �  J5  Z5  �  �3  �3   +pop_back ,_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv �5  �5  �   ,!  E_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ 8�  6  )6  �  �  �  ,�   ,!  [_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_yy 8�  �6  �6  �  �  �  ,�  �  �   ,!  t_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy 8�  7  7  �  �  �  �  �   ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc 8�  u7  �7  �  �  �  �      �   ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc 8�  �7  �7  �  �  �  �  �    ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ 8�  �8  �8  �  �3  �3  ,�   ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y 8�  9  39  �  �3  �3  �  �   ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ 8�  �9  �9  �  �3  �3  �   ,!  �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc 8�  K:  e:  �  �3  �3  �  �    ,!  /_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ 8�  �:  ;  �  �3  �3  �  �   ,!  :_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ 8��        �;  �;  �  �3  �3  �  �   ,!  E_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ 8�  0<  J<  �  �3  �3  �  �   ,!  P_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ 8�  �<  �<  �  �3  �3  r  r   ,!  i_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE 8�  =  �=  �  r  r  g   %_M_replace_aux �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc 8�  �=  >  �  �  �  �  �    %_M_replace �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replaceEyyPKcy 8�  ~>  �>  �  �  �  �  �   %_M_append �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy 8�  �>  ?  �  �  �   -copy �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy �  `?  u?  �  �  �  �   �      +swap �_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ �?  �?  �  8�   -c_str �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5c_strEv �  *@  0@  �   -data �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv �  �@  �@  �   -get_allocator �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv Q  �@  �@  �   ,  	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy �  QA  fA  �  �  �  �   ,  	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERKS4_y �  �A  �A  �  ,�  �   ,  <	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy �  &B  6B  �  �  �   ,  M	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy �  �B  �B  �  �   �   ,�  Z	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y �  �B  C  �  ,�  �   ,�  |	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy �  ^C  sC  �  �  �  �      �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy �  �C  �C  �  �  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy �  1D  AD  �  �   �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y �  �D  �D  �  ,�  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcyy �  E  +E  �  �  �  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy �  �E  �E  �  �  �   ,�  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEcy �  �E  F  �  �   �   ,(  �	_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y �  mF  }F  �  ,�  �   ,(   
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy �  �F  �F  �  �  �  �   ,(  .
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcy �  SG  cG  �  �  �   ,(�        B
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy �  �G  �G  �  �   �   ,�  P
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofERKS4_y �  8H  HH  �  ,�  �   ,�  s
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy �  �H  �H  �  �  �  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy �  (I  8I  �  �  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy �  �I  �I  �  �   �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y �  J  !J  �  ,�  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy �  �J  �J  �  �  �  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy �  �J  K  �  �  �   ,�  �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not�      _ofEcy �  qK  �K  �  �   �   -substr �
_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy   �K  �K  �  �  �   ,_  _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ l  FL  QL  �  ,�   ,_  e_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ l  �L  �L  �  �  �  ,�   ,_  _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy l  "M  AM  �  �  �  ,�  �  �   ,_  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEPKc l  �M  �M  �  �   ,_  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc l   N  N  �  �  �  �   ,_  �_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKcy l  qN  �N  �  �  �  �  �   /�  �   0  NY  0�  �a     string J!   1
A	  2@��  2�1  2���  2�։  2���  2��  2�9�  2�^�  2�|�  2���  2���  2�؊  2��  2��  2�I�  2�j�  2���  2���  �      2�֋  2��  2��  2�4�  2�T�  2�{�  2���  2���  2��  2��  2�-�  2�M�  2�r�  2���  2���  2�͍  2��  2�
�  2�;�  2�T�  2�x�  2���  2���  2��  2��  2�?�  2�g�  2���  2���  2�Ώ  2��  2��  2�0�  2�U�  2�{�  2���  2���  2�א  2���  2��  2�3�  2�Q�  3v�  3	��  3
ʑ  3?�  3{�  3�  3!-�  3%v�  3&��  3'ʑ  �  V
4Q  4�  Y_ZNSt9nothrow_tC4Ev -Q  �    �P  5nothrow ]_ZSt7nothrow 4Q  6__exception_ptr 	4�U  7�  	O�U  _M_exception_object 	Q��   8�  	S_ZNSt15__exception_ptr13exception_ptrC4EPv �Q  �Q  ��  ��    _M_addref 	U_ZNSt15__exception_ptr13exception_ptr9_M_addrefEv &R  ,R  ��    _M_release 	V_ZNSt15__exception_ptr13exception_ptr10_M_releaseEv wR  }R  ��   !_M_get 	X_ZNKSt15__exception_ptr13exception_ptr6_M_getEv ��  �R  �R  ��   9�  	`_ZNSt15__exception_ptr13exception_ptrC4Ev S  S  ��   9�  	b_ZNSt15__exception_ptr13exception_ptrC4ERKS0_ JS  US  ���        �   9�  	e_ZNSt15__exception_ptr13exception_ptrC4EDn �S  �S  ��  IV   9�  	i_ZNSt15__exception_ptr13exception_ptrC4EOS0_ �S  �S  ��  �   :|  	v_ZNSt15__exception_ptr13exception_ptraSERKS0_ #�  (T  3T  ��  �   :|  	z_ZNSt15__exception_ptr13exception_ptraSEOS0_ #�  uT  �T  ��  �   ;~exception_ptr 	�_ZNSt15__exception_ptr13exception_ptrD4Ev �T  �T  ��  l   ;swap 	�_ZNSt15__exception_ptr13exception_ptr4swapERS0_ U  U  ��  #�   <operator bool 	�_ZNKSt15__exception_ptr13exception_ptrcvbEv )�  iU  oU  ��   =__cxa_exception_type 	�_ZNKSt15__exception_ptr13exception_ptr20__cxa_exception_typeEv 6�  �U  ��    nQ  2	I�U   2	9nQ  >rethrow_exception 	E_ZSt17rethrow_exceptionNSt15__exception_ptr13exception_ptrE IV  nQ   nullptr_t 
�
�  ?type_info [V  integral_constant<bool, false> E6W  @value G-1�  A  H-)�  !operator std::integral_constant<bool, false>::value_type J_ZNKSt17integral_constantIbLb0EEcvbEv �V  W  "W  <�   B_Tp )�  C__v )�    kV  integral_�      constant<bool, true> EX  @value G-1�  A  H-)�  !operator std::integral_constant<bool, true>::value_type J_ZNKSt17integral_constantIbLb1EEcvbEv pW  �W  �W  B�   B_Tp )�  C__v )�   ;W  D__swappable_details u	__is_integer<long double> dX  E�  �ZX  F8    B_Tp ��   __is_integer<double> �X  E�  ��X  F8    B_Tp /�   __is_integer<float> �X  E�  ��X  F8    B_Tp ^�   �  L
Y  4�  L+_ZNSt21piecewise_construct_tC4Ev Y  W�    �X  Gpiecewise_construct O5Y   H__debug 2char_traits<char> ]  '  _ZNSt11char_traitsIcE6assignERcRKc �Y  �  ��   I^  !�   �Y  (eq  _ZNSt11char_traitsIcE2eqERKcS2_ )�  �Y  ��  ��   (lt $_ZNSt11char_traitsIcE2ltERKcS2_ )�  -Z  ��  ��   J_  ,_ZNSt11char_traitsIcE7compareEPKcS2_y l  tZ  ��  ��  ]   Jh  :_ZNSt11char_traitsIcE6lengthEPKc ]  �Z  ��   J  D_ZNSt11char_traitsIcE4findEPKcyRS1_ ��  �Z  ��  ]  ��   (move R_ZNSt11char_traitsIcE4moveEPcPKcy ��  5[  ��  ��  ]   (copy Z�      _ZNSt11char_traitsIcE4copyEPcPKcy ��  y[  ��  ��  ]   J  b_ZNSt11char_traitsIcE6assignEPcyc ��  �[  ��  ]  �Y   Jo  j_ZNSt11char_traitsIcE12to_char_typeERKi �Y  �[  ��   It  !l  �[  J�  p_ZNSt11char_traitsIcE11to_int_typeERKc �[  K\  ��   J�  t_ZNSt11char_traitsIcE11eq_int_typeERKiS2_ )�  �\  ��  ��   Keof x_ZNSt11char_traitsIcE3eofEv �[  (not_eof |_ZNSt11char_traitsIcE7not_eofERKi �[  �\  ��   /�  �    size_t 
��   char_traits<wchar_t> ��`  '  �_ZNSt11char_traitsIwE6assignERwRKw j]  ��  ��   I^  �!�  j]  (eq �_ZNSt11char_traitsIwE2eqERKwS2_ )�  �]  ��  ��   (lt �_ZNSt11char_traitsIwE2ltERKwS2_ )�  �]  ��  ��   J_  �_ZNSt11char_traitsIwE7compareEPKwS2_y l  9^  ��  ��  ]   Jh  �_ZNSt11char_traitsIwE6lengthEPKw ]  q^  ��   J  �_ZNSt11char_traitsIwE4findEPKwyRS1_ ��  �^  ��  ]  ��   (move �_ZNSt11char_traitsIwE4moveEPwPKwy ��  �^  ��  ��  ]   (copy �_ZNSt11char_traitsIwE4copyEPwPKwy ��  >_  ��  ��      �  ]   J  �_ZNSt11char_traitsIwE6assignEPwyw ��  �_  ��  ]  j]   Jo  �_ZNSt11char_traitsIwE12to_char_typeERKt j]  �_  ��   It  �!1  �_  J�  �_ZNSt11char_traitsIwE11to_int_typeERKw �_  `  ��   J�  �_ZNSt11char_traitsIwE11eq_int_typeERKtS2_ )�  V`  ��  ��   Keof �_ZNSt11char_traitsIwE3eofEv �_  (not_eof �_ZNSt11char_traitsIwE7not_eofERKt �_  �`  ��   /�  �   20��  21ڒ  22��  23�  25�  26�  27C�  28n�  2:=�  2;h�  2<��  2=  2?��  2@  2Bʒ  2C�  2D�  2E,�  2G�  2H-�  2IX�  2J��  2LR�  2M~�  2N��  2Oؓ  2Q��  2R  25  26�  27	�  ptrdiff_t 
��   allocator<char> lmb  L�n   9@  �_ZNSaIcEC4Ev b  b  ��   9@  �_ZNSaIcEC4ERKS_ 5b  @b  ��  ��   M~allocator �_ZNSaIcED4Ei ab  ��  l    �a  2ז  2��  2��  2���  2��  2�+�  2�C�  2���  2���  2�  2�ߙ  2���  2�#�  2�G�  2�k�  2�y�  2���  2���  2�њ  2���  2��  2�5�  2���  2��      .r  2�T�  2�r�  2�֛  2���  2���  2���  2b��  2cԔ  2e�  2f-�  2gG�  2h_�  2iy�  2j��  2k��  2lҜ  2m��  2n�  2q4�  2r\�  2s��  2t��  2uĝ  2v�  2x�  2y�  2|,�  2~D�  2Z�  2�u�  2���  2���  2�  2�ܞ  2���  2�!�  2�B�  2�b�  2�s�  2���  2���  2�ҟ  2��  2��  2�?�  2�d�  2���  2���  allocator_traits<std::allocator<char> > �g  I�  ��  J�  �_ZNSt16allocator_traitsISaIcEE8allocateERS0_y �d  ;e  Ԡ  Me   I  �,�a  ;e  I  �$]  J�  �_ZNSt16allocator_traitsISaIcEE8allocateERS0_yPKv �d  �e  Ԡ  Me  �e   const_void_pointer �-z�  '5  �_ZNSt16allocator_traitsISaIcEE10deallocateERS0_Pcy f  Ԡ  �d  Me   J�  �_ZNSt16allocator_traitsISaIcEE8max_sizeERKS0_ Me  ]f  ڠ   (select_on_container_copy_construction �_ZNSt16allocator_traitsISaIcEE37select_on_container_copy_constructionERKS0_ ;e  �f  ڠ   I  ��   I�  �'�  rebind_alloc �%�a  /�  �a   initiali�      zer_list<char> /�h  �  6�  _M_array :<g     5]  _M_len ;[g  �  >_ZNSt16initializer_listIcEC4EPKcy �g  �g  >�  �g  [g   )  7�  9�  B_ZNSt16initializer_listIcEC4Ev �g  �g  >�   Nsize G_ZNKSt16initializer_listIcE4sizeEv [g  6h  <h  D�   Nbegin K_ZNKSt16initializer_listIcE5beginEv �g  wh  }h  D�   Nend O_ZNKSt16initializer_listIcE3endEv �g  �h  �h  D�   B_E �    g  ?reverse_iterator<__gnu_cxx::__normal_iterator<char*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > > ?reverse_iterator<__gnu_cxx::__normal_iterator<char const*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > > O_V2 GPG�i  Qios_base �j  RInit [+Init __ZNSt8ios_base4InitC4Ev 7j  =j  J�   +~Init `_ZNSt8ios_base4InitD4Ev ij  tj  J�  l   S_S_refcount ce�  S_S_synced_with_stdio d)�    2RP�  2S[  2T1  2\b�  2e��  2h��  2i��  Qbasic_ostream<char, std::char_traits<char> > &k  /�  �   0�        NY   Qbasic_ostream<wchar_t, std::char_traits<wchar_t> > qk  /�  �  0  ]   Qbasic_istream<char, std::char_traits<char> > �k  /�  �   0  NY   Qbasic_istream<wchar_t, std::char_traits<wchar_t> > l  /�  �  0  ]   istream �!qk  5cin <_ZSt3cin l  ostream �!�j  5cout =_ZSt4cout &l  5cerr >_ZSt4cerr &l  5clog ?_ZSt4clog &l  wistream �#�k  5wcin B_ZSt4wcin {l  wostream �#&k  5wcout C_ZSt5wcout �l  5wcerr D_ZSt5wcerr �l  5wclog E_ZSt5wclog �l  T__ioinit J j  Uabs N_ZSt3abse ��  0m  ��   Uabs J_ZSt3absf ^�  Pm  ^�   Uabs F_ZSt3absd /�  pm  /�   Uabs =_ZSt3absx �   �m  �    Uabs 8_ZSt3absl x  �m  x   Udiv �_ZSt3divll �  �m  x  x   iterator_traits<char*> �$n  A�  �+�a  A�  �+�  AO  �+��  /g  �   Viterator_traits<char const*> �A�  �+�a  A�  �+�  AO  �+��  /g  �    W__gnu_cxx 
��  X__cxx11 
A1
A�n  2�v�  3��  3ʑ  H__ops #2,]  2-�a  new_allocator<char> :�q  9�  O_ZN9__gnu_cxx13new_allocatorIc�      EC4Ev $o  *o  ��   9�  Q_ZN9__gnu_cxx13new_allocatorIcEC4ERKS1_ co  no  ��  ��   ;~new_allocator V_ZN9__gnu_cxx13new_allocatorIcED4Ev �o  �o  ��  l   �  ?�  Naddress Y_ZNK9__gnu_cxx13new_allocatorIcE7addressERc �o  p  p  ��  p   O  A��  �  @�  Naddress ]_ZNK9__gnu_cxx13new_allocatorIcE7addressERKc #p  vp  �p  ��  �p   d  B��  :�  c_ZN9__gnu_cxx13new_allocatorIcE8allocateEyPKv �o  �p  �p  ��  �p  z�     =]  95  t_ZN9__gnu_cxx13new_allocatorIcE10deallocateEPcy /q  ?q  ��  �o  �p   :�  �_ZNK9__gnu_cxx13new_allocatorIcE8max_sizeEv �p  �q  �q  ��   B_Tp �    �n  __numeric_traits_integer<int> 7�q  Y�  :s  Y1  ;s  Y�  ?1�  Y  @s  /X  l   2���  2�T�  2�r�  2���  2���  2�֛  2���  Udiv �_ZN9__gnu_cxx3divExx ��  ^r  �   �    2��  2�?�  2�d�  2���  2���  __alloc_traits<std::allocator<char>, char>  2
�u  2 2
Ze  2 2
�d  2 2
�e  2 2
f  �d   U_S_select_on_copy  ^_ZN9__gnu_cxx14__alloc_�      traitsISaIcEcE17_S_select_on_copyERKS1_ �a  Cs  ��   Z_S_on_swap  a_ZN9__gnu_cxx14__alloc_traitsISaIcEcE10_S_on_swapERS1_S3_ �s  �  �   [_S_propagate_on_copy_assign  d_ZN9__gnu_cxx14__alloc_traitsISaIcEcE27_S_propagate_on_copy_assignEv )�  [_S_propagate_on_move_assign  g_ZN9__gnu_cxx14__alloc_traitsISaIcEcE27_S_propagate_on_move_assignEv )�  [_S_propagate_on_swap  j_ZN9__gnu_cxx14__alloc_traitsISaIcEcE20_S_propagate_on_swapEv )�  [_S_always_equal  m_ZN9__gnu_cxx14__alloc_traitsISaIcEcE15_S_always_equalEv )�  [_S_nothrow_move  p_ZN9__gnu_cxx14__alloc_traitsISaIcEcE15_S_nothrow_moveEv )�  A   :5�f  ju  A�   ;5�d  A�   <5�f  A   =5Me  AO   @5�  Ad   A5�  rebind<char>  t�u  other  uA�f  B_Tp �    /�  �a   \__normal_iterator<char*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > !�|}  ]  !��   )�  !_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4Ev �v  �v  s�   *�  !_ZN9__gnu_cxx17__nor�      mal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4ERKS1_ [w  fw  s�  y�   ^O  !2n  ,@  !_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEdeEv fw  �w  �w  �   ^�  !2n  ,�  !_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEptEv �w  px  vx  �   ,�  !!_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEv ��  �x  �x  s�   ,�  !(_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEi �u  by  my  s�  l   ,�  !-_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEv ��  �y  �y  s�   ,�  !4_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEi �u  Yz  dz  s�  l   ,�  !9_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEixEx fw  �z  �z  �  �z   ^�  !8�m  ,  !=_ZN�      9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEpLEx ��  d{  o{  s�  �z   ,J  !A_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEplEx �u  �{  �{  �  �z   ,�  !E_ZN9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmIEx ��  a|  l|  s�  �z   ,T  !I_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmiEx �u  �|  �|  �  �z   -base !M_ZNK9__gnu_cxx17__normal_iteratorIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEE4baseEv y�  c}  i}  �   /g  �  /D     �u  \__normal_iterator<char const*, std::__cxx11::basic_string<char, std::char_traits<char>, std::allocator<char> > > !�"�  ]  !��   )�  !_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4Ev {~  �~  [�   *�  !_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEC4ERKS2_ �~     �      [�  a�   ^O  !2^n  ,@  !_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEdeEv    �  �  g�   ^�  !2Rn  ,�  !_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEptEv �  �  �  g�   ,�  !!_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEv m�  ��  ��  [�   ,�  !(_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEppEi �}   �  �  [�  l   ,�  !-_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEv m�  �  ��  [�   ,�  !4_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmmEi �}  ��  �  [�  l   ,�  !9_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEixEx    y�  ��  g�  ��   ^�  !8Fn  ,  !=_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcES�      aIcEEEEpLEx m�  �  �  [�  ��   ,J  !A_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEplEx �}  ��  ��  g�  ��   ,�  !E_ZN9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmIEx m�  �  �  [�  ��   ,T  !I_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEmiEx �}  ��  ��  g�  ��   -base !M_ZNK9__gnu_cxx17__normal_iteratorIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEE4baseEv a�  	�  �  g�   /g  �  /D     �}  __numeric_traits_floating<float> d��  Y  gs  Y�  j1�  YY  ks  Y�  ls  /X  ^�   __numeric_traits_floating<double> d��  Y  gs  Y�  j1�  YY  ks  Y�  ls  /X  /�   __numeric_traits_floating<long double> dZ�  Y  gs  Y�  j1�  YY  ks  Y�  ls  /X  ��   __numeric_traits_integer<long unsigned int> 7Ɇ  Y�  :�  Y1  ;�  Y�  ?1�  Y  @s  /X  �   __numeric_traits_integer<ch�      ar> 7+�  Y�  :�   Y1  ;�   Y�  ?1�  Y  @s  /X  �    __numeric_traits_integer<short int> 7��  Y�  :�  Y1  ;�  Y�  ?1�  Y  @s  /X  ��   V__numeric_traits_integer<long long int> 7Y�  :	  Y1  ;	  Y�  ?1�  Y  @s  /X  �     _iobuf 0")
��  _ptr "*�   _cnt "+	l  _base ",�  _flag "-	l  _file ".	l  _charbuf "/	l   _bufsiz "0	l  $_tmpfname "1�  ( FILE "3��  ___imp__pctype "���  �  ___imp__wctype "���  ___imp__pwctype "���  short int ��  tm $"Q
��  
tm_sec "R	l   
tm_min "S	l  
tm_hour "T	l  
tm_mday "U	l  
tm_mon "V	l  
tm_year "W	l  
tm_wday "X	l  
tm_yday "Y	l  
tm_isdst "Z	l    �  mbstate_t "�l  ��  `btowc "�1  ։  l   `fgetwc "1  ��  ��   ��  `fgetws "�  �  �  l  ��   `fputwc "1  9�  �  ��   `fputws "l  X�  X�  ��   �  `fwide "�l  |�  ��  l   afwprintf "Il  ��  ��  X�  b afwscanf "%l  ��  ��  X�  b `getwc "1  ؊  ��   cgetw�      char "1  `mbrlen "��   �  �  �   �   �   �  ��  `mbrtowc "��   I�  �  �  �   �   `mbsinit "�l  d�  d�   ��  `mbsrtowcs "��   ��  �  ��  �   �   �  `putwc "	1  ��  �  ��   `putwchar "
1  ֋  �   d}  #>l  �  �  X�  b d}  #"l  �  �  �   X�  b aswscanf "l  4�  X�  X�  b `ungetwc "1  T�  1  ��   avfwprintf "_l  {�  ��  X�  �    avfwscanf "?l  ��  ��  X�  �    d  #3l  ��  �  X�  �    d  #l  �  �  �   X�  �    avswscanf "1l  �  X�  X�  �    avwprintf "fl  -�  X�  �    avwscanf "8l  M�  X�  �    `wcrtomb "��   r�  �  �  �   ewcscat $��  ��  �  X�   ewcscmp $�l  ��  X�  X�   ewcscoll $�l  ͍  X�  X�   ewcscpy $��  �  �  X�   ewcscspn $��   
�  X�  X�   `wcsftime "e�   5�  �  �   X�  5�   ��  ewcslen $��   T�  X�   ewcsncat $��  x�  �  X�  �    ewcsncmp $�l  ��  X�  X�  �    ewcsncpy $��  ��  �  X�  �    `wcsrtombs "��   쎜        �  �  �   �   X�  ewcsspn $��   �  X�  X�   awcstod "�/�  /�  X�  9�   double �  awcstof "�^�  ^�  X�  9�   float ewcstok $��  ��  �  X�   `wcstol "�x  ��  X�  9�  l   `wcstoul "��  Ώ  X�  9�  l   ewcsxfrm $��   �  �  X�  �    `wctob "�l  �  1   `wmemcmp "�l  0�  X�  X�  �    `wmemcpy "��  U�  �  X�  �    `wmemmove "��  {�  �  X�  �    `wmemset "��  ��  �  �  �    awprintf "Tl  ��  X�  b awscanf "l  א  X�  b ewcschr $�"�  ��  X�  �   ewcspbrk $�"�  �  X�  X�   ewcsrchr $�"�  3�  X�  �   ewcsstr $�"�  Q�  X�  X�   `wmemchr "�"�  v�  X�  �  �    `wcstold "���  ��  X�  9�   long double `wcstoll "�'�   ʑ  X�  9�  l   `wcstoull "�0�   �  X�  9�  l   �P  fnQ  �U  g�U  hdecltype(nullptr) inQ  gnQ  bool )�  fV  6W  X  signed char �X  j$Y  6__gnu_debug 8�  P:BY   g�Y  g�Y  �Y  �Y  g\  gj]  gw]  w]  j]  g�_  int8_t %#H�  ui�      nt8_t %$�  int16_t %%��  uint16_t %&@  int32_t %'l  uint32_t %(�  int64_t %)&�   uint64_t %*0�   int_least8_t %-H�  uint_least8_t %.�  int_least16_t %/��  uint_least16_t %0@  int_least32_t %1l  uint_least32_t %2�  int_least64_t %3&�   uint_least64_t %40�   int_fast8_t %:H�  uint_fast8_t %;�  int_fast16_t %<��  uint_fast16_t %=@  int_fast32_t %>l  uint_fast32_t %?�  int_fast64_t %@&�   uint_fast64_t %A0�   intmax_t %D&�   uintmax_t %E0�   char16_t char32_t fpos_t &h%�   Ԕ  esetlocale P�  	�  l  �   klocaleconv Q!�  �  '�  l ___newclmap 'P�  ___newcumap 'Q�  ___ptlocinfo 'R�  ___ptmbcinfo 'S�  ___globallocalestatus 'Tl  ___locale_changed 'Ul  ___initiallocinfo 'V(�  ___initiallocalestructinfo 'W  ___imp___mb_cur_max '��  �  m�  n�  l   ___security_cookie (}  n>�  ��   3�  o_pthread_key_dest )#_�  >�  _Atomic_word * l  ��  p�n  g�q  �q  g�   g�   �a  gmb  _div_t +;ז  quot +<	l�         rem +=	l   div_t +>��  _ldiv_t +@�  quot +A
x   rem +B
x   ldiv_t +C�  �  1�  �     __sys_errlist +�&!�  __sys_nerr +�$l  o__imp___argc +�  o__imp___argv +��  ��  �  o__imp___wargv +!��  9�  o__imp__environ +'��  o__imp__wenviron +,��  o__imp__pgmptr +2��  o__imp__wpgmptr +79�  o__imp__osplatform +<(�  �  o__imp__osver +A(�  o__imp__winver +F(�  o__imp__winmajor +K(�  o__imp__winminor +P(�  q+�7lldiv_t ��  
quot +�0�    
rem +�6�    lldiv_t +�=��  __amblksiz ,5�  `atexit +�l  ��  �   `atof +�/�  �  �   `atoi +�l  +�  �   `atol +�x  C�  �   `bsearch +���  r�  z�  z�  �   �   r�   x�  rl  ��  z�  z�   `div +�ז  ��  l  l   `getenv +��    �   `ldiv +��  ߙ  x  x   `mblen +�l  ��  �  �    `mbstowcs +��   #�  �  �  �    `mbtowc +�l  G�  �  �  �    sqsort +�k�  ��  �   �   r�   crand +�l  ssrand +���  �   astrtod +� /�  ��  �  ��   `strtol +�x  �      њ  �  ��  l   `strtoul +��  ��  �  ��  l   esystem (Ul  �  �   `wcstombs +��   5�  �  X�  �    `wctomb +�l  T�  �  �   `lldiv +�%��  r�  �   �    `atoll +�(�   ��  �   `strtoll +�(�   ��  �  ��  l   `strtoull +�1�   ֛  �  ��  l   astrtof +�^�  ��  �  ��   `strtold +�'��  �  �  ��   sclearerr &B-�  ��   `fclose &Cl  G�  ��   `feof &Jl  _�  ��   `ferror &Kl  y�  ��   `fflush &Ll  ��  ��   `fgetc &Ml  ��  ��   `fgetpos &Ol  ̜  ��  ̜   Ԕ  `fgets &Q�  ��  �  l  ��   `fopen &X��  �  �  �   afprintf &Nl  4�  ��  �  b `fread &]�   \�  ��  �   �   ��   `freopen &^��  ��  �  �  ��   afscanf &!l  ��  ��  �  b `fseek &al  ĝ  ��  x  l   `fsetpos &_l  �  ��  �   �  `ftell &bx  �  ��   `getc &�l  �  ��   cgetchar &�l  `gets &��  D�  �   sperror &�Z�  �   aprintf &Yl  u�  �  b eremove -�l  ��  �   erename -�l  ��  �  �   srewind &�      �  ��   ascanf &l  ܞ  �  b ssetbuf &���  ��  �   `setvbuf &�l  !�  ��  �  l  �    asprintf &dl  B�  �  �  b asscanf &l  b�  �  �  b ctmpfile &���  `tmpnam &��  ��  �   `ungetc &�l  ��  l  ��   avfprintf &ol  ҟ  ��  �  �    avprintf &vl  �  �  �    avsprintf &}l  �  �  �  �    asnprintf &�l  ?�  �  �   �  b avfscanf &@l  d�  ��  �  �    avscanf &9l  ��  �  �    avsnprintf &�l  ��  �  �   �  �    avsscanf &2l  Ԡ  �  �  �    g;e  gHe  g�a  gju  gvu  e  i�a  �   �  �      �N  g�  gQ  g^  g�N  i  g  g  �h   j  wctrans_t .��  `iswctype "#l  ��  1  [   etowctrans .�1  ��  1  P�   ewctrans .�P�  ��  �   ewctype .�[  ס  �   t�l  	@�L     _PHNDLR /?�  _XCPT_ACTION /A
B�  XcptNum /B�   SigNum /C	l  XcptAction /D�   ��  M�  l __XcptActTab /GB�  __XcptActTabCount /Hl  __XcptActTabSize /Il  __First_FPE_Indx /Jl  __N�      um_FPE /Kl  DWORD 0��  _GUID 1�  Data1 1�   Data2 1@  Data3 1@  Data4 1�   �  %�  �    GUID 1ɢ  %�  IID 1S%�  7�  CLSID 1[%�  H�  FMTID 1b%�  [�  oGUID_MAX_POWER_SAVINGS 2�2�  oGUID_MIN_POWER_SAVINGS 2�2�  oGUID_TYPICAL_POWER_SAVINGS 2�2�  oNO_SUBGROUP_GUID 2�2�  oALL_POWERSCHEMES_GUID 2�2�  oGUID_POWERSCHEME_PERSONALITY 2�2�  oGUID_ACTIVE_POWERSCHEME 2�2�  oGUID_IDLE_RESILIENCY_SUBGROUP 2�2�  oGUID_IDLE_RESILIENCY_PERIOD 2�2�  oGUID_DISK_COALESCING_POWERDOWN_TIMEOUT 2�2�  oGUID_EXECUTION_REQUIRED_REQUEST_TIMEOUT 2�2�  oGUID_VIDEO_SUBGROUP 2�2�  oGUID_VIDEO_POWERDOWN_TIMEOUT 2�2�  oGUID_VIDEO_ANNOYANCE_TIMEOUT 2�2�  oGUID_VIDEO_ADAPTIVE_PERCENT_INCREASE 2�2�  oGUID_VIDEO_DIM_TIMEOUT 2�2�  oGUID_VIDEO_ADAPTIVE_POWERDOWN 2�2�  oGUID_MONITOR_POWER_ON 2�2�  oGUID_DEVICE_POWER_POLICY_VIDEO_BRIGHTNESS 2�2�  oGUID_DEVICE_POWER_POLICY_VIDEO_DIM_BRIGHTNESS 2�2�  oGUID_VIDEO_CURRENT_MONITOR_BRIGHTNESS 2�2�  oGUID_VIDEO_ADAP�      TIVE_DISPLAY_BRIGHTNESS 2�2�  oGUID_CONSOLE_DISPLAY_STATE 2�2�  oGUID_ALLOW_DISPLAY_REQUIRED 2�2�  oGUID_VIDEO_CONSOLE_LOCK_TIMEOUT 2�2�  oGUID_ADAPTIVE_POWER_BEHAVIOR_SUBGROUP 2�2�  oGUID_NON_ADAPTIVE_INPUT_TIMEOUT 2�2�  oGUID_DISK_SUBGROUP 2�2�  oGUID_DISK_POWERDOWN_TIMEOUT 2�2�  oGUID_DISK_IDLE_TIMEOUT 2�2�  oGUID_DISK_BURST_IGNORE_THRESHOLD 2�2�  oGUID_DISK_ADAPTIVE_POWERDOWN 2�2�  oGUID_SLEEP_SUBGROUP 2�2�  oGUID_SLEEP_IDLE_THRESHOLD 2�2�  oGUID_STANDBY_TIMEOUT 2�2�  oGUID_UNATTEND_SLEEP_TIMEOUT 2�2�  oGUID_HIBERNATE_TIMEOUT 2�2�  oGUID_HIBERNATE_FASTS4_POLICY 2�2�  oGUID_CRITICAL_POWER_TRANSITION 2�2�  oGUID_SYSTEM_AWAYMODE 2�2�  oGUID_ALLOW_AWAYMODE 2�2�  oGUID_ALLOW_STANDBY_STATES 2�2�  oGUID_ALLOW_RTC_WAKE 2�2�  oGUID_ALLOW_SYSTEM_REQUIRED 2�2�  oGUID_SYSTEM_BUTTON_SUBGROUP 2�2�  oGUID_POWERBUTTON_ACTION 2�2�  oGUID_SLEEPBUTTON_ACTION 2�2�  oGUID_USERINTERFACEBUTTON_ACTION 2�2�  oGUID_LIDCLOSE_ACTION 2�2�  oGUID_LIDOPEN_POWERSTATE 2�2��        oGUID_BATTERY_SUBGROUP 2�2�  oGUID_BATTERY_DISCHARGE_ACTION_0 2�2�  oGUID_BATTERY_DISCHARGE_LEVEL_0 2�2�  oGUID_BATTERY_DISCHARGE_FLAGS_0 2�2�  oGUID_BATTERY_DISCHARGE_ACTION_1 2�2�  oGUID_BATTERY_DISCHARGE_LEVEL_1 2�2�  oGUID_BATTERY_DISCHARGE_FLAGS_1 2�2�  oGUID_BATTERY_DISCHARGE_ACTION_2 2�2�  oGUID_BATTERY_DISCHARGE_LEVEL_2 2�2�  oGUID_BATTERY_DISCHARGE_FLAGS_2 2�2�  oGUID_BATTERY_DISCHARGE_ACTION_3 2�2�  oGUID_BATTERY_DISCHARGE_LEVEL_3 2�2�  oGUID_BATTERY_DISCHARGE_FLAGS_3 2�2�  oGUID_PROCESSOR_SETTINGS_SUBGROUP 2�2�  oGUID_PROCESSOR_THROTTLE_POLICY 2�2�  oGUID_PROCESSOR_THROTTLE_MAXIMUM 2�2�  oGUID_PROCESSOR_THROTTLE_MINIMUM 2�2�  oGUID_PROCESSOR_ALLOW_THROTTLING 2�2�  oGUID_PROCESSOR_IDLESTATE_POLICY 2�2�  oGUID_PROCESSOR_PERFSTATE_POLICY 2�2�  oGUID_PROCESSOR_PERF_INCREASE_THRESHOLD 2�2�  oGUID_PROCESSOR_PERF_DECREASE_THRESHOLD 2�2�  oGUID_PROCESSOR_PERF_INCREASE_POLICY 2�2�  oGUID_PROCESSOR_PERF_DECREASE_POLICY 2�2�  oGUID_PROCESSOR_PERF_INCRE�      ASE_TIME 2�2�  oGUID_PROCESSOR_PERF_DECREASE_TIME 2�2�  oGUID_PROCESSOR_PERF_TIME_CHECK 2�2�  oGUID_PROCESSOR_PERF_BOOST_POLICY 2�2�  oGUID_PROCESSOR_PERF_BOOST_MODE 2�2�  oGUID_PROCESSOR_IDLE_ALLOW_SCALING 2�2�  oGUID_PROCESSOR_IDLE_DISABLE 2�2�  oGUID_PROCESSOR_IDLE_STATE_MAXIMUM 2�2�  oGUID_PROCESSOR_IDLE_TIME_CHECK 2�2�  oGUID_PROCESSOR_IDLE_DEMOTE_THRESHOLD 2�2�  oGUID_PROCESSOR_IDLE_PROMOTE_THRESHOLD 2�2�  oGUID_PROCESSOR_CORE_PARKING_INCREASE_THRESHOLD 2�2�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_THRESHOLD 2�2�  oGUID_PROCESSOR_CORE_PARKING_INCREASE_POLICY 2 2�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_POLICY 22�  oGUID_PROCESSOR_CORE_PARKING_MAX_CORES 22�  oGUID_PROCESSOR_CORE_PARKING_MIN_CORES 22�  oGUID_PROCESSOR_CORE_PARKING_INCREASE_TIME 22�  oGUID_PROCESSOR_CORE_PARKING_DECREASE_TIME 22�  oGUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_DECREASE_FACTOR 22�  oGUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_THRESHOLD 22�  oGUID_PROCESSOR_CORE_PARKING_A�      FFINITY_WEIGHTING 22�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_DECREASE_FACTOR 2	2�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_THRESHOLD 2
2�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_WEIGHTING 22�  oGUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_THRESHOLD 22�  oGUID_PROCESSOR_PARKING_CORE_OVERRIDE 22�  oGUID_PROCESSOR_PARKING_PERF_STATE 22�  oGUID_PROCESSOR_PARKING_CONCURRENCY_THRESHOLD 22�  oGUID_PROCESSOR_PARKING_HEADROOM_THRESHOLD 22�  oGUID_PROCESSOR_PERF_HISTORY 22�  oGUID_PROCESSOR_PERF_LATENCY_HINT 22�  oGUID_PROCESSOR_DISTRIBUTE_UTILITY 22�  oGUID_SYSTEM_COOLING_POLICY 22�  oGUID_LOCK_CONSOLE_ON_WAKE 22�  oGUID_DEVICE_IDLE_POLICY 22�  oGUID_ACDC_POWER_SOURCE 22�  oGUID_LIDSWITCH_STATE_CHANGE 22�  oGUID_BATTERY_PERCENTAGE_REMAINING 22�  oGUID_GLOBAL_USER_PRESENCE 22�  oGUID_SESSION_DISPLAY_STATUS 22�  oGUID_SESSION_USER_PRESENCE 22�  oGUID_IDLE_BACKGROUND_TASK 22�  oGUID_BACKGROUND_TASK_NOTIFICATION 2�      2�  oGUID_APPLAUNCH_BUTTON 22�  oGUID_PCIEXPRESS_SETTINGS_SUBGROUP 2 2�  oGUID_PCIEXPRESS_ASPM_POLICY 2!2�  oGUID_ENABLE_SWITCH_FORCED_SHUTDOWN 2"2�  oPPM_PERFSTATE_CHANGE_GUID 2 2�  oPPM_PERFSTATE_DOMAIN_CHANGE_GUID 2!2�  oPPM_IDLESTATE_CHANGE_GUID 2"2�  oPPM_PERFSTATES_DATA_GUID 2#2�  oPPM_IDLESTATES_DATA_GUID 2$2�  oPPM_IDLE_ACCOUNTING_GUID 2%2�  oPPM_IDLE_ACCOUNTING_EX_GUID 2&2�  oPPM_THERMALCONSTRAINT_GUID 2'2�  oPPM_PERFMON_PERFSTATE_GUID 2(2�  oPPM_THERMAL_POLICY_CHANGE_GUID 2)2�  RPC_IF_HANDLE 3B��  24'�  243ז  244�  `abs +l  ָ  l   246��  246m  2460m  246Pm  246pm  246�m  247��  248�  249+�  24:C�  24<.r  24<��  24<�m  24>��  24@  24Cߙ  24D��  24E#�  24GG�  24Hk�  24Jy�  24K��  24L��  24Mњ  24N��  24P�  24Q5�  _IWinTypesBase_v0_1_c_ifspec 5)��  _IWinTypesBase_v0_1_s_ifspec 5*��  _IID_IUnknown 6=C�  _IID_AsyncIUnknown 6�2�  oIID_IClassFactory 6m2�  oIID_IMarshal 7n2�  oIID_INoMarshal 7U2�  oIID_IAgileObje�      ct 7�2�  oIID_IAgileReference 7�2�  oIID_IMarshal2 7-2�  oIID_IMalloc 7�2�  oIID_IStdMarshalInfo 7i2�  oIID_IExternalConnection 7�2�  oIID_IMultiQI 7G2�  oIID_AsyncIMultiQI 7�2�  oIID_IInternalUnknown 72�  oIID_IEnumUnknown 7h2�  oIID_IEnumString 72�  oIID_ISequentialStream 7�2�  oIID_IStream 7M2�  oIID_IRpcChannelBuffer 7�	2�  oIID_IRpcChannelBuffer2 7;
2�  oIID_IAsyncRpcChannelBuffer 7�
2�  oIID_IRpcChannelBuffer3 72�  oIID_IRpcSyntaxNegotiate 7�2�  oIID_IRpcProxyBuffer 7�2�  oIID_IRpcStubBuffer 7V2�  oIID_IPSFactoryBuffer 72�  oIID_IChannelHook 7�2�  oIID_IClientSecurity 7�2�  oIID_IServerSecurity 7m2�  oIID_IRpcOptions 72�  oIID_IGlobalOptions 7�2�  oIID_ISurrogate 7!2�  oIID_IGlobalInterfaceTable 7�2�  oIID_ISynchronize 72�  oIID_ISynchronizeHandle 7�2�  oIID_ISynchronizeEvent 7�2�  oIID_ISynchronizeContainer 7A2�  oIID_ISynchronizeMutex 7�2�  oIID_ICancelMethodCalls 72�  oIID_IAsyncManager 7�2�  oIID_ICallFactory 72�  o�      IID_IRpcHelper 7f2�  oIID_IReleaseMarshalBuffers 7�2�  oIID_IWaitMultiple 7,2�  oIID_IAddrTrackingControl 7�2�  oIID_IAddrExclusionControl 7�2�  oIID_IPipeByte 7h2�  oIID_IPipeLong 7�2�  oIID_IPipeDouble 7J2�  oIID_IComThreadingInfo 7$2�  oIID_IProcessInitControl 7�2�  oIID_IFastRundown 72�  oIID_IMarshalingStream 7J2�  oIID_ICallbackWithNoReentrancyToApplicationSTA 7	2�  _GUID_NULL 8C�  _CATID_MARSHALER 8C�  _IID_IRpcChannel 8C�  _IID_IRpcStub 8C�  _IID_IStubManager 8C�  _IID_IRpcProxy 8C�  _IID_IProxyManager 8C�  _IID_IPSFactory 8C�  _IID_IInternalMoniker 8C�  _IID_IDfReserved1 8C�  _IID_IDfReserved2 8C�  _IID_IDfReserved3 8C�  _CLSID_StdMarshal 8V�  _CLSID_AggStdMarshal 8V�  _CLSID_StdAsyncActManager 8V�  _IID_IStub 8C�  _IID_IProxy 8C�  _IID_IEnumGeneric 8C�  _IID_IEnumHolder 8C�  _IID_IEnumCallback 8 C�  _IID_IOleManager 8!C�  _IID_IOlePresObj 8"C�  _IID_IDebug 8#C�  _IID_IDebugStream 8$C�  _CLSID_PSGenObject 8%V�  _CLSID_PSCl�      ientSite 8&V�  _CLSID_PSClassObject 8'V�  _CLSID_PSInPlaceActive 8(V�  _CLSID_PSInPlaceFrame 8)V�  _CLSID_PSDragDrop 8*V�  _CLSID_PSBindCtx 8+V�  _CLSID_PSEnumerators 8,V�  _CLSID_StaticMetafile 8-V�  _CLSID_StaticDib 8.V�  _CID_CDfsVolume 8/V�  _CLSID_DCOMAccessControl 80V�  _CLSID_GlobalOptions 81V�  _CLSID_StdGlobalInterfaceTable 82V�  _CLSID_ComBinding 83V�  _CLSID_StdEvent 84V�  _CLSID_ManualResetEvent 85V�  _CLSID_SynchronizeContainer 86V�  _CLSID_AddrControl 87V�  _CLSID_CCDFormKrnl 88V�  _CLSID_CCDPropertyPage 89V�  _CLSID_CCDFormDialog 8:V�  _CLSID_CCDCommandButton 8;V�  _CLSID_CCDComboBox 8<V�  _CLSID_CCDTextBox 8=V�  _CLSID_CCDCheckBox 8>V�  _CLSID_CCDLabel 8?V�  _CLSID_CCDOptionButton 8@V�  _CLSID_CCDListBox 8AV�  _CLSID_CCDScrollBar 8BV�  _CLSID_CCDGroupBox 8CV�  _CLSID_CCDGeneralPropertyPage 8DV�  _CLSID_CCDGenericPropertyPage 8EV�  _CLSID_CCDFontPropertyPage 8FV�  _CLSID_CCDColorPropertyPage 8GV�  _CLSID_CCDLabelPropertyPage 8HV�  _CLSID_CCDCheckBoxPro�      pertyPage 8IV�  _CLSID_CCDTextBoxPropertyPage 8JV�  _CLSID_CCDOptionButtonPropertyPage 8KV�  _CLSID_CCDListBoxPropertyPage 8LV�  _CLSID_CCDCommandButtonPropertyPage 8MV�  _CLSID_CCDComboBoxPropertyPage 8NV�  _CLSID_CCDScrollBarPropertyPage 8OV�  _CLSID_CCDGroupBoxPropertyPage 8PV�  _CLSID_CCDXObjectPropertyPage 8QV�  _CLSID_CStdPropertyFrame 8RV�  _CLSID_CFormPropertyPage 8SV�  _CLSID_CGridPropertyPage 8TV�  _CLSID_CWSJArticlePage 8UV�  _CLSID_CSystemPage 8VV�  _CLSID_IdentityUnmarshal 8WV�  _CLSID_InProcFreeMarshaler 8XV�  _CLSID_Picture_Metafile 8YV�  _CLSID_Picture_EnhMetafile 8ZV�  _CLSID_Picture_Dib 8[V�  _GUID_TRISTATE 8\2�  _IWinTypes_v0_1_c_ifspec 9(��  _IWinTypes_v0_1_s_ifspec 9)��  oIID_IMallocSpy :�2�  oIID_IBindCtx ::2�  oIID_IEnumMoniker :J 2�  oIID_IRunnableObject :� 2�  oIID_IRunningObjectTable :�!2�  oIID_IPersist :i"2�  oIID_IPersistStream :�"2�  oIID_IMoniker :j#2�  oIID_IROTData :X%2�  oIID_IEnumSTATSTG :�%2�  oIID_IStorage :X&2�  oIID_IPersistFile�       :A(2�  oIID_IPersistStorage :�(2�  oIID_ILockBytes :�)2�  oIID_IEnumFORMATETC :�*2�  oIID_IEnumSTATDATA :l+2�  oIID_IRootStorage :,2�  oIID_IAdviseSink :�,2�  oIID_AsyncIAdviseSink :s-2�  oIID_IAdviseSink2 :�.2�  oIID_AsyncIAdviseSink2 :./2�  oIID_IDataObject :�/2�  oIID_IDataAdviseHolder :12�  oIID_IMessageFilter :�12�  oFMTID_SummaryInformation :]2i�  oFMTID_DocSummaryInformation :_2i�  oFMTID_UserDefinedProperties :a2i�  oFMTID_DiscardableInformation :c2i�  oFMTID_ImageSummaryInformation :e2i�  oFMTID_AudioSummaryInformation :g2i�  oFMTID_VideoSummaryInformation :i2i�  oFMTID_MediaFileSummaryInformation :k2i�  oIID_IClassActivator :s22�  oIID_IFillLockBytes :�22�  oIID_IProgressNotify :�32�  oIID_ILayoutStorage :�32�  oIID_IBlockingLock :�42�  oIID_ITimeAndNoticeControl :�42�  oIID_IOplockStorage :N52�  oIID_IDirectWriterLock :�52�  oIID_IUrlMon :M62�  oIID_IForegroundTransfer :�62�  oIID_IThumbnailExtractor :72�  oIID_IDummyHICONIncluder :�72�  oIID_IProcessLoc�      k :�72�  oIID_ISurrogateService :H82�  oIID_IInitializeSpy :�82�  oIID_IApartmentShutdown :�92�  _IID_IOleAdviseHolder ;�2�  oIID_IOleCache ;b2�  oIID_IOleCache2 ;)2�  oIID_IOleCacheControl ;�2�  oIID_IParseDisplayName ;<2�  oIID_IOleContainer ;�2�  oIID_IOleClientSite ;2�  oIID_IOleObject ;�2�  oIOLETypes_v0_0_c_ifspec ;���  oIOLETypes_v0_0_s_ifspec ;���  oIID_IOleWindow ;$2�  oIID_IOleLink ;�2�  oIID_IOleItemContainer ;�2�  oIID_IOleInPlaceUIWindow ;v	2�  oIID_IOleInPlaceActiveObject ;
2�  oIID_IOleInPlaceFrame ;�
2�  oIID_IOleInPlaceObject ;�2�  oIID_IOleInPlaceSite ;�2�  oIID_IContinue ;�2�  oIID_IViewObject ;�2�  oIID_IViewObject2 ;*2�  oIID_IDropSource ;�2�  oIID_IDropTarget ;[2�  oIID_IDropSourceNotify ;�2�  oIID_IEnumOLEVERB ;v2�  _IID_IServiceProvider <9C�  _IOleAutomationTypes_v1_0_c_ifspec =���  _IOleAutomationTypes_v1_0_s_ifspec =���  oIID_ICreateTypeInfo =;2�  oIID_ICreateTypeInfo2 =b2�  oIID_ICreateTypeLib =�2�  oIID_ICreateTyp�      eLib2 =�2�  oIID_IDispatch =�	2�  oIID_IEnumVARIANT =�
2�  oIID_ITypeComp =52�  oIID_ITypeInfo =�2�  oIID_ITypeInfo2 =P2�  oIID_ITypeLib =�2�  oIID_ITypeLib2 ==2�  oIID_ITypeChangeEvents =a2�  oIID_IErrorInfo =�2�  oIID_ICreateErrorInfo =}2�  oIID_ISupportErrorInfo = 2�  oIID_ITypeFactory =u2�  oIID_ITypeMarshal =�2�  oIID_IRecordInfo =�2�  oIID_IErrorLog = 2�  oIID_IPropertyBag =z2�  ___MIDL_itf_msxml_0000_v0_0_c_ifspec >���  ___MIDL_itf_msxml_0000_v0_0_s_ifspec >���  _LIBID_MSXML >�C�  oIID_IXMLDOMImplementation > C�  oIID_IXMLDOMNode >'C�  oIID_IXMLDOMDocumentFragment >�C�  oIID_IXMLDOMDocument >fC�  oIID_IXMLDOMNodeList >uC�  oIID_IXMLDOMNamedNodeMap >�C�  oIID_IXMLDOMCharacterData >C�  oIID_IXMLDOMAttribute >�C�  oIID_IXMLDOMElement >C�  oIID_IXMLDOMText >�C�  oIID_IXMLDOMComment >%C�  oIID_IXMLDOMProcessingInstruction >�C�  oIID_IXMLDOMCDATASection >C�  oIID_IXMLDOMDocumentType >�C�  oIID_IXMLDOMNotation >C�  oIID_IXMLDOMEntity�       >C�  oIID_IXMLDOMEntityReference >�C�  oIID_IXMLDOMParseError >a	C�  oIID_IXTLRuntime >�	C�  oDIID_XMLDOMDocumentEvents >=
C�  oCLSID_DOMDocument >\
V�  oCLSID_DOMFreeThreadedDocument >`
V�  oIID_IXMLHttpRequest >g
C�  oCLSID_XMLHTTPRequest >�
V�  oIID_IXMLDSOControl >�
C�  oCLSID_XMLDSOControl >V�  oIID_IXMLElementCollection >C�  oIID_IXMLDocument >JC�  oIID_IXMLDocument2 >�C�  oIID_IXMLElement >$C�  oIID_IXMLElement2 >�C�  oIID_IXMLAttribute >�C�  oIID_IXMLError >C�  oCLSID_XMLDocument >.V�  oCLSID_SBS_StdURLMoniker ?~C�  oCLSID_SBS_HttpProtocol ?C�  oCLSID_SBS_FtpProtocol ?�C�  oCLSID_SBS_GopherProtocol ?�C�  oCLSID_SBS_HttpSProtocol ?�C�  oCLSID_SBS_FileProtocol ?�C�  oCLSID_SBS_MkProtocol ?�C�  oCLSID_SBS_UrlMkBindCtx ?�C�  oCLSID_SBS_SoftDistExt ?�C�  oCLSID_SBS_CdlProtocol ?�C�  oCLSID_SBS_ClassInstallFilter ?�C�  oCLSID_SBS_InternetSecurityManager ?�C�  oCLSID_SBS_InternetZoneManager ?�C�  oIID_IAsyncMoniker ?�C�  oCLSID_StdURLMon�      iker ?�C�  oCLSID_HttpProtocol ?�C�  oCLSID_FtpProtocol ?�C�  oCLSID_GopherProtocol ?�C�  oCLSID_HttpSProtocol ?�C�  oCLSID_FileProtocol ?�C�  oCLSID_MkProtocol ?�C�  oCLSID_StdURLProtocol ?�C�  oCLSID_UrlMkBindCtx ?�C�  oCLSID_CdlProtocol ?�C�  oCLSID_ClassInstallFilter ?�C�  oIID_IAsyncBindCtx ?�C�  oIID_IPersistMoniker ?P2�  oIID_IMonikerProp ?!2�  oIID_IBindProtocol ?2�  oIID_IBinding ?�2�  oIID_IBindStatusCallback ?u2�  oIID_IBindStatusCallbackEx ?�2�  oIID_IAuthenticate ?d2�  oIID_IAuthenticateEx ?�2�  oIID_IHttpNegotiate ?A2�  oIID_IHttpNegotiate2 ?�2�  oIID_IHttpNegotiate3 ?;	2�  oIID_IWinInetFileStream ?�	2�  oIID_IWindowForBindingUI ?0
2�  oIID_ICodeInstall ?�
2�  oIID_IWinInetInfo ?�2�  oIID_IHttpSecurity ?2�  oIID_IWinInetHttpInfo ?y2�  oIID_IWinInetHttpTimeouts ?�2�  oSID_BindHost ?52�  oIID_IBindHost ??2�  oIID_IInternet ?M2�  oIID_IInternetBindInfo ?�2�  oIID_IInternetBindInfoEx ?&2�  oIID_IInternetProtocolRoot ?�2�  �      oIID_IInternetProtocol ?�2�  oIID_IInternetProtocolSink ?2�  oIID_IInternetProtocolSinkStackable ?�2�  oIID_IInternetSession ??2�  oIID_IInternetThreadSwitch ?H2�  oIID_IInternetPriority ?�2�  oIID_IInternetProtocolInfo ?N2�  oCLSID_InternetSecurityManager ?�C�  oCLSID_InternetZoneManager ?�C�  oIID_IInternetSecurityMgrSite ?�2�  oIID_IInternetSecurityManager ?i2�  oIID_IInternetHostSecurityManager ?!2�  oIID_IInternetZoneManager ?�"2�  oCLSID_SoftDistExt ?�&C�  oIID_ISoftDistExt ?�&2�  oIID_ICatalogFileInfo ?x'2�  oIID_IDataFilter ?�'2�  oIID_IEncodingFilterFactory ?�(2�  oGUID_CUSTOM_CONFIRMOBJECTSAFETY ?3)2�  oIID_IWrappedProtocol ?A)2�  oIID_IGetBindHandle ?�)2�  oIID_IBindCallbackRedirect ?*2�  oIID_IPropertyStorage @�2�  oIID_IPropertySetStorage @2�  oIID_IEnumSTATPROPSTG @�2�  oIID_IEnumSTATPROPSETSTG @D2�  _IID_StdOle AC�  _GUID_DEVINTERFACE_DISK B2�  _GUID_DEVINTERFACE_CDROM B2�  _GUID_DEVINTERFACE_PARTITION B2�  _GUID_DEVINTERFACE_TAPE B�      2�  _GUID_DEVINTERFACE_WRITEONCEDISK B2�  _GUID_DEVINTERFACE_VOLUME B2�  _GUID_DEVINTERFACE_MEDIUMCHANGER B2�  _GUID_DEVINTERFACE_FLOPPY B2�  _GUID_DEVINTERFACE_CDCHANGER B2�  _GUID_DEVINTERFACE_STORAGEPORT B2�  _GUID_DEVINTERFACE_COMPORT B2�  _GUID_DEVINTERFACE_SERENUM_BUS_ENUMERATOR B2�  _SCARD_IO_REQUEST C���  dwProtocol C���   cbPciLength C���   SCARD_IO_REQUEST C�`�  ��  _g_rgSCardT0Pci D%.��  _g_rgSCardT1Pci D%=��  _g_rgSCardRawPci D%L��  _IID_IPrintDialogCallback E2�  _IID_IPrintDialogServices E2�  2F�N  2F6l  �}  g�  "�  g�}  �u  g�  |}  g�u  u_ZNSt17integral_constantIbLb0EE5valueE �V   u_ZNSt17integral_constantIbLb1EE5valueE bW  v_ZN9__gnu_cxx24__numeric_traits_integerIiE5__minE �q  ����xw_ZN9__gnu_cxx24__numeric_traits_integerIiE5__maxE �q  ���u_ZN9__gnu_cxx25__numeric_traits_floatingIfE16__max_exponent10E u�  &x_ZN9__gnu_cxx25__numeric_traits_floatingIdE16__max_exponent10E څ  4x_ZN9__gnu_cxx25__numeric_traits_floatingIeE16__max_exponent10�      E D�  Du_ZN9__gnu_cxx24__numeric_traits_integerImE8__digitsE ��   u_ZN9__gnu_cxx24__numeric_traits_integerIcE5__maxE ��  v_ZN9__gnu_cxx24__numeric_traits_integerIsE5__minE X�  ��~x_ZN9__gnu_cxx24__numeric_traits_integerIsE5__maxE d�  �v_ZN9__gnu_cxx24__numeric_traits_integerIxE5__minE ��  ���������y_ZN9__gnu_cxx24__numeric_traits_integerIxE5__maxE ˇ  �������z_GLOBAL__sub_I_disk.cpp g@            �{__static_initialization_and_destruction_0 +@     <       �0�  |__initialize_p l  � |__priority l  � z__tcf_0 @            � *         �@     R�@       S  �  ��     GNU C17 8.1.0 -mtune=core2 -march=nocona -g -g -g -O2 -O2 -O2 -fno-ident -fbuilding-libgcc -fno-stack-protector ../../../../../src/gcc-8.1.0/libgcc/libgcc2.c C:\mingw810\x86_64-810-posix-seh-rt_v6-rev0\build\gcc-8.1.0\x86_64-w64-mingw32\libgcc �  char   long long unsigned int long long int uintptr_t K,  wchar_t b_  short unsigned int int u  long int   O  u  u�      nsigned int long unsigned int unsigned char long double double float __imp___mb_cur_max s�    �  )  	    _sys_errlist �&  _sys_nerr �$u  
__imp___argc �  
__imp___argv |  �  �  
__imp___wargv !�  �  �  
__imp__environ '|  
__imp__wenviron ,�  
__imp__pgmptr 2�  
__imp__wpgmptr 7�  
__imp__osplatform <&  �  
__imp__osver A&  
__imp__winver F&  
__imp__winmajor K&  
__imp__winminor P&  _amblksiz 5�  __security_cookie }=  optarg #�  optind 1u  opterr 6u  optopt :u    �  _daylight zu  _dstbias {�  _timezone |�  �  C  	   _tzname }3  
daylight u  
timezone �  
tzname 3  short int hashval_t *�  htab_hash /�  �  �  �  �   �  htab_eq 6�  �  u  �  �  �   htab_hash_pointer ��  htab_eq_pointer ��  stringop_alg �  
�  no_stringop  libcall rep_prefix_1_byte rep_prefix_4_byte rep_prefix_8_by�      te loop_1_byte loop unrolled_loop vector_loop last_alg 	 0  �  �   �  
unspec_strings X�  
unspecv_strings ��  stringop_strategy 	�k  max 	�|   alg 	��  noalign 	�	u   $  stringop_algs 4	��  unknown_size 	��   size 	��   k  �  	   �  processor_costs �	��  add 	�|   lea 	�|  shift_var 	�|  shift_const 	�|  mult_init 	��  mult_bit 	�|  $divide 	��  (movsx 	�u  <movzx 	�u  @large_insn 	�|  Dmove_ratio 	�|  Hmovzbl_load 	�|  Lint_load 	�  Pint_store 	�  \fp_move 	�|  hfp_load 	�  lfp_store 	�  xmmx_move 	 |  �mmx_load 	  �mmx_store 	  �xmm_move 	|  �ymm_move 	|  �zmm_move 	|  �sse_load 	�  �sse_unaligned_load 		�  �sse_store 	
�  �sse_unaligned_store 	�  �mmxsse_to_integer 	|  �ssemmx_to_integer 	|  �gather_static 	|  �gather_per_elt 	|   scatter_static 	|  scatter_per_elt 	|  l1_cache_size 	|  �      l2_cache_size 	|  prefetch_block 	|  simultaneous_prefetches 	|  branch_cost 	|  fadd 	|   fmul 	|  $fdiv 	|  (fabs 	|  ,fchs 	|  0fsqrt 	|  4sse_op 	"|  8addss 	#|  <mulss 	$|  @mulsd 	%|  Dfmass 	&|  Hfmasd 	'|  Ldivss 	(|  Pdivsd 	)|  Tsqrtss 	*|  Xsqrtsd 	+|  \reassoc_int 	,|  `reassoc_fp 	,|  dreassoc_vec_int 	,&|  hreassoc_vec_fp 	,7|  lmemcpy 	3!  pmemset 	3"!  xcond_taken_branch_cost 	4|  �cond_not_taken_branch_cost 	6|  � �  |  �  	   �  |    	   �  |    	     p  
ix86_cost 	:&:  �  
ix86_size_cost 	;%�  ix86_tune_indices �  	�z  X86_TUNE_SCHEDULE  X86_TUNE_PARTIAL_REG_DEPENDENCY X86_TUNE_SSE_PARTIAL_REG_DEPENDENCY X86_TUNE_SSE_SPLIT_REGS X86_TUNE_PARTIAL_FLAG_REG_STALL X86_TUNE_MOVX X86_TUNE_MEMORY_MISMATCH_STALL X86_TUNE_FUSE_CMP_AND_BRANCH_32 X86_TUNE_FUSE_CMP_AND_BRANCH_64 X86_�      TUNE_FUSE_CMP_AND_BRANCH_SOFLAGS 	X86_TUNE_FUSE_ALU_AND_BRANCH 
X86_TUNE_ACCUMULATE_OUTGOING_ARGS X86_TUNE_PROLOGUE_USING_MOVE X86_TUNE_EPILOGUE_USING_MOVE X86_TUNE_USE_LEAVE X86_TUNE_PUSH_MEMORY X86_TUNE_SINGLE_PUSH X86_TUNE_DOUBLE_PUSH X86_TUNE_SINGLE_POP X86_TUNE_DOUBLE_POP X86_TUNE_PAD_SHORT_FUNCTION X86_TUNE_PAD_RETURNS X86_TUNE_FOUR_JUMP_LIMIT X86_TUNE_SOFTWARE_PREFETCHING_BENEFICIAL X86_TUNE_LCP_STALL X86_TUNE_READ_MODIFY X86_TUNE_USE_INCDEC X86_TUNE_INTEGER_DFMODE_MOVES X86_TUNE_OPT_AGU X86_TUNE_AVOID_LEA_FOR_ADDR X86_TUNE_SLOW_IMUL_IMM32_MEM X86_TUNE_SLOW_IMUL_IMM8 X86_TUNE_AVOID_MEM_OPND_FOR_CMOVE  X86_TUNE_SINGLE_STRINGOP !X86_TUNE_MISALIGNED_MOVE_STRING_PRO_EPILOGUES "X86_TUNE_USE_SAHF #X86_TUNE_USE_CLTD $X86_TUNE_USE_BT %X86_TUNE_AVOID_FALSE_DEP_FOR_BMI &X86_TUNE_ADJUST_UNROLL 'X86_TUNE_ONE_IF_CONV_INSN (X86_TUNE_USE_HIMODE_FIOP )X86_TUNE_USE_SIMODE_FIOP *X86_TUNE_USE_FFREEP +X86_TUNE_EXT_80387_CONSTANTS ,X86_TUNE_GENERAL_REGS_SSE_S�      PILL -X86_TUNE_SSE_UNALIGNED_LOAD_OPTIMAL .X86_TUNE_SSE_UNALIGNED_STORE_OPTIMAL /X86_TUNE_SSE_PACKED_SINGLE_INSN_OPTIMAL 0X86_TUNE_SSE_TYPELESS_STORES 1X86_TUNE_SSE_LOAD0_BY_PXOR 2X86_TUNE_INTER_UNIT_MOVES_TO_VEC 3X86_TUNE_INTER_UNIT_MOVES_FROM_VEC 4X86_TUNE_INTER_UNIT_CONVERSIONS 5X86_TUNE_SPLIT_MEM_OPND_FOR_FP_CONVERTS 6X86_TUNE_USE_VECTOR_FP_CONVERTS 7X86_TUNE_USE_VECTOR_CONVERTS 8X86_TUNE_SLOW_PSHUFB 9X86_TUNE_AVOID_4BYTE_PREFIXES :X86_TUNE_USE_GATHER ;X86_TUNE_AVOID_128FMA_CHAINS <X86_TUNE_AVX256_UNALIGNED_LOAD_OPTIMAL =X86_TUNE_AVX256_UNALIGNED_STORE_OPTIMAL >X86_TUNE_AVX128_OPTIMAL ?X86_TUNE_AVX256_OPTIMAL @X86_TUNE_DOUBLE_WITH_ADD AX86_TUNE_ALWAYS_FANCY_MATH_387 BX86_TUNE_UNROLL_STRLEN CX86_TUNE_SHIFT1 DX86_TUNE_ZERO_EXTEND_WITH_AND EX86_TUNE_PROMOTE_HIMODE_IMUL FX86_TUNE_FAST_PREFIX GX86_TUNE_READ_MODIFY_WRITE HX86_TUNE_MOVE_M1_VIA_OR IX86_TUNE_NOT_UNPAIRABLE JX86_TUNE_PARTIAL_REG_STALL KX86_TUNE_PROMOTE_QIMODE LX86_TUNE_PROMOTE_HI_REGS MX86_TUNE_HIMODE_MATH N�      X86_TUNE_SPLIT_LONG_MOVES OX86_TUNE_USE_XCHGB PX86_TUNE_USE_MOV0 QX86_TUNE_NOT_VECTORMODE RX86_TUNE_AVOID_VECTOR_DECODE SX86_TUNE_BRANCH_PREDICTION_HINTS TX86_TUNE_QIMODE_MATH UX86_TUNE_PROMOTE_QI_REGS VX86_TUNE_EMIT_VZEROUPPER WX86_TUNE_LAST X �  �  	  W 
ix86_tune_features 	�z  ix86_arch_indices �  	"1  X86_ARCH_CMOV  X86_ARCH_CMPXCHG X86_ARCH_CMPXCHG8B X86_ARCH_XADD X86_ARCH_BSWAP X86_ARCH_LAST  �  A  	   
ix86_arch_features 	,1  
x86_prefetch_sse 	;�  _dont_use_tree_here_ 
x86_mfence 	Y�  w  reg_class �  	*�  NO_REGS  AREG DREG CREG BREG SIREG DIREG AD_REGS CLOBBERED_REGS Q_REGS 	NON_Q_REGS 
TLS_GOTBASE_REGS INDEX_REGS LEGACY_REGS GENERAL_REGS FP_TOP_REG FP_SECOND_REG FLOAT_REGS SSE_FIRST_REG NO_REX_SSE_REGS SSE_REGS EVEX_SSE_REGS BND_REGS ALL_SSE_REGS MMX_REGS FP_TOP_SSE_REGS FP_SECOND_SSE_REGS FLOAT_SSE_REGS FLOAT_INT_REGS INT_SSE_REGS FLOAT_INT_SSE_REGS MASK_EVEX_REGS MASK�      _REGS  MOD4_SSE_REGS !ALL_REGS "LIM_REG_CLASSES # �  |  �  	  P �  
dbx_register_map 	=�  
dbx64_register_map 	>�  
svr4_dbx_register_map 	?�  processor_type �  	��  PROCESSOR_GENERIC  PROCESSOR_I386 PROCESSOR_I486 PROCESSOR_PENTIUM PROCESSOR_LAKEMONT PROCESSOR_PENTIUMPRO PROCESSOR_PENTIUM4 PROCESSOR_NOCONA PROCESSOR_CORE2 PROCESSOR_NEHALEM 	PROCESSOR_SANDYBRIDGE 
PROCESSOR_HASWELL PROCESSOR_BONNELL PROCESSOR_SILVERMONT PROCESSOR_KNL PROCESSOR_KNM PROCESSOR_SKYLAKE PROCESSOR_SKYLAKE_AVX512 PROCESSOR_CANNONLAKE PROCESSOR_ICELAKE_CLIENT PROCESSOR_ICELAKE_SERVER PROCESSOR_INTEL PROCESSOR_GEODE PROCESSOR_K6 PROCESSOR_ATHLON PROCESSOR_K8 PROCESSOR_AMDFAM10 PROCESSOR_BDVER1 PROCESSOR_BDVER2 PROCESSOR_BDVER3 PROCESSOR_BDVER4 PROCESSOR_BTVER1 PROCESSOR_BTVER2  PROCESSOR_ZNVER1 !PROCESSOR_max " 
ix86_tune 		  
ix86_arch 		  
ix86_preferred_stack_boundary 			�  
ix86_incoming_stack_boundary 	
	�  �  o  	�        P _  
regclass_map 		o  signed char UQItype {�  �  __int128 __int128 unsigned complex float complex double  complex long double _Float128  complex _Float128 �  ;  	  � +  
__popcount_tab �;  
__clz_tab ;  func_ptr *  k  �   __CTOR_LIST__ /|  __DTOR_LIST__ 0|  �  9	
	 J     �  :	
	xJ      7s   O  GNU C17 8.1.0 -mtune=core2 -march=nocona -g -g -g -O2 -O2 -O2 -fno-ident -fbuilding-libgcc -fno-stack-protector -fexceptions ../../../../../src/gcc-8.1.0/libgcc/unwind-seh.c C:\mingw810\x86_64-810-posix-seh-rt_v6-rev0\build\gcc-8.1.0\x86_64-w64-mingw32\libgcc `�@     '      5  char %  long long unsigned int long long int uintptr_t K,2  wchar_t b  short unsigned int   int �  long int pthreadlocinfo �(�  �  threadlocaleinfostruct `�z  C  ��   	lc_codepage ��  	lc_collate_cp ��  	lc_handle ��  	lc_id �	�  $	lc_category �  H
lc_clike ��  
mb_cur_max �      ��  
lconv_intl_refcount ��  
lconv_num_refcount ��  
lconv_mon_refcount ��   
lconv �#  (
ctype1_refcount ��  0
ctype1 �)  8
pctype �/  @
pclmap �5  H
pcumap �5  P
lc_time_curr �a  X pthreadmbcinfo �%�  �  threadmbcinfostruct localeinfo_struct ��  	locinfo ��   	mbcinfo �z   _locale_tstruct ��  tagLC_ID �V  	wLanguage �   	wCountry �  	wCodePage �   LC_ID �   ��  	locale ��   	wlocale ��  C  �
�  	wrefcount �
�   %  o  �  unsigned int �  �  2   long unsigned int V    2   e    2   lconv     �  L  unsigned char ;  __lc_time_data Q  long double double float __imp___mb_cur_max s�  �  �  2    _sys_errlist �&�  _sys_nerr �$�  __imp___argc �  __imp___argv     �  __imp___wargv !*  0  �  __imp__environ '  __imp__wenviron ,*  __imp__pgmptr 2  __�      imp__wpgmptr 70  __imp__osplatform <�  �  __imp__osver A�  __imp__winver F�  __imp__winmajor K�  __imp__winminor P�  _amblksiz 5�  .  9  �   __security_cookie }]  optarg #�  optind 1�  opterr 6�  optopt :�  -  �  _daylight z�  _dstbias {�  _timezone |�  �  �  2   _tzname }�  daylight �  timezone �  tzname �  short int hashval_t *�  htab_hash /T  Z  0  i  i   o  htab_eq 6�  �  �  �  i  i   htab_hash_pointer �B  htab_eq_pointer �p  stringop_alg �  |	  no_stringop  libcall rep_prefix_1_byte rep_prefix_4_byte rep_prefix_8_byte loop_1_byte loop unrolled_loop vector_loop last_alg 	 �  �  �	   �	  unspec_strings 	X�	  unspecv_strings 	��	  stringop_strategy 
�	
  max 
��   alg 
�|	  noalign 
�	�   �	  stringop_algs 4
�J
  unknown_size 
�|	   size 
�Z
   	
  Z
  2   J
  processor_costs �
�{  �      add 
��   lea 
��  shift_var 
��  shift_const 
��  mult_init 
��  mult_bit 
��  $divide 
��  (movsx 
��  <movzx 
��  @large_insn 
��  Dmove_ratio 
��  Hmovzbl_load 
��  Lint_load 
��  Pint_store 
��  \fp_move 
��  hfp_load 
��  lfp_store 
��  x	mmx_move 
 �  �	mmx_load 
�  �	mmx_store 
�  �	xmm_move 
�  �	ymm_move 
�  �	zmm_move 
�  �	sse_load 
�  �	sse_unaligned_load 
	�  �	sse_store 

�  �	sse_unaligned_store 
�  �	mmxsse_to_integer 
�  �	ssemmx_to_integer 
�  �	gather_static 
�  �
gather_per_elt 
�   
scatter_static 
�  
scatter_per_elt 
�  
l1_cache_size 
�  
l2_cache_size 
�  
prefetch_block 
�  
simultaneous_prefetches 
�  
branch_cost 
�  
fadd 
�   
fmul 
�  $
fdiv 
�  (
fabs 
�  ,
fchs 
�  0
fsqrt 
�  4
sse_op 
"�  8
addss 
#�  <
mulss 
$�  @
mulsd 
%�  D
fmass 
&�  H
fmasd 
'�  L
divss 
(�      �  P
divsd 
)�  T
sqrtss 
*�  X
sqrtsd 
+�  \
reassoc_int 
,�  `
reassoc_fp 
,�  d
reassoc_vec_int 
,&�  h
reassoc_vec_fp 
,7�  l
memcpy 
3�  p
memset 
3"�  x
cond_taken_branch_cost 
4�  �
cond_not_taken_branch_cost 
6�  � _
  �  �  2   �  �  �  2   �  �  �  2   �  
  ix86_cost 
:&�  {  ix86_size_cost 
;%{  ;    2  W ix86_tune_features 
��  ;  2  2   ix86_arch_features 
,"  x86_prefetch_sse 
;;  _dont_use_tree_here_ x86_mfence 
Y�  h  reg_class �  
*�  NO_REGS  AREG DREG CREG BREG SIREG DIREG AD_REGS CLOBBERED_REGS Q_REGS 	NON_Q_REGS 
TLS_GOTBASE_REGS INDEX_REGS LEGACY_REGS GENERAL_REGS FP_TOP_REG FP_SECOND_REG FLOAT_REGS SSE_FIRST_REG NO_REX_SSE_REGS SSE_REGS EVEX_SSE_REGS BND_REGS ALL_SSE_REGS MMX_REGS FP_TOP_SSE_REGS FP_SECOND_SSE_REGS FLOAT_SSE_REGS FLOAT_INT_REGS INT_SSE_REGS FLOAT_INT_SSE_REGS MASK_EVEX_REGS MASK_REGS�        MOD4_SSE_REGS !ALL_REGS "LIM_REG_CLASSES # �  �  �  2  P �  dbx_register_map 
=�  dbx64_register_map 
>�  svr4_dbx_register_map 
?�  processor_type �  
��  PROCESSOR_GENERIC  PROCESSOR_I386 PROCESSOR_I486 PROCESSOR_PENTIUM PROCESSOR_LAKEMONT PROCESSOR_PENTIUMPRO PROCESSOR_PENTIUM4 PROCESSOR_NOCONA PROCESSOR_CORE2 PROCESSOR_NEHALEM 	PROCESSOR_SANDYBRIDGE 
PROCESSOR_HASWELL PROCESSOR_BONNELL PROCESSOR_SILVERMONT PROCESSOR_KNL PROCESSOR_KNM PROCESSOR_SKYLAKE PROCESSOR_SKYLAKE_AVX512 PROCESSOR_CANNONLAKE PROCESSOR_ICELAKE_CLIENT PROCESSOR_ICELAKE_SERVER PROCESSOR_INTEL PROCESSOR_GEODE PROCESSOR_K6 PROCESSOR_ATHLON PROCESSOR_K8 PROCESSOR_AMDFAM10 PROCESSOR_BDVER1 PROCESSOR_BDVER2 PROCESSOR_BDVER3 PROCESSOR_BDVER4 PROCESSOR_BTVER1 PROCESSOR_BTVER2  PROCESSOR_ZNVER1 !PROCESSOR_max " ix86_tune 
	  ix86_arch 
	  ix86_preferred_stack_boundary 
		�  ix86_incoming_stack_boundary 

	�  �  `  2  P �      P  regclass_map 
	`  _PHNDLR ?(  _XCPT_ACTION A
�  XcptNum B�   SigNum C	�  XcptAction D{   �  �   _XcptActTab G�  _XcptActTabCount H�  _XcptActTabSize I�  _First_FPE_Indx J�  _Num_FPE K�  V  _EXCEPTION_RECORD ��
  	ExceptionCode �
m   	ExceptionFlags �
m  	ExceptionRecord �
!P  	ExceptionAddress �
�  	NumberParameters �
m  	ExceptionInformation �
F"      _CONTEXT ��%7  	P1Home ��   	P2Home ��  	P3Home ��  	P4Home ��  	P5Home ��   	P6Home ��  (	ContextFlags �m  0	MxCsr �m  4	SegCs �
`  8	SegDs �
`  :	SegEs �
`  <	SegFs �
`  >	SegGs �
`  @	SegSs �
`  B	EFlags �m  D	Dr0 ��  H	Dr1 ��  P	Dr2 ��  X	Dr3 ��  `	Dr6 ��  h	Dr7 ��  p	Rax ��  x	Rcx ��  �	Rdx ��  �	Rbx ��  �	Rsp ��  �	Rbp ��  �	Rsi ��  �	Rdi ��  �	R8 ��  �	R9 ��  �	R10 ��  �	R11 ��  �	R12 ��  �	R13 ��  �	R14 ��  �	R15 ��      �  �	Rip ��  � Y!   !VectorRegister ��!   
VectorControl ��  �
DebugControl ��  �
LastBranchToRip ��  �
LastBranchFromRip ��  �
LastExceptionToRip ��  �
LastExceptionFromRip ��  � ULONG �  UCHAR ;  BYTE �;  WORD �  DWORD ��  __imp__pctype +�  )  __imp__wctype ;�  __imp__pwctype G�  L  �   �  __newclmap P�  __newcumap Q�  __ptlocinfo R�  __ptmbcinfo Sz  __globallocalestatus T�  __locale_changed U�  __initiallocinfo V(�  __initiallocalestructinfo W�  signed char ULONG_PTR 1.2  ULONG64 �.2  DWORD64 �.2  PVOID �  LONGLONG �%L  ULONGLONG �.2  _GUID T  Data1 �   Data2   Data3   Data4 T   ;  d  2   GUID   d  IID Sd  v  CLSID [d  �  FMTID bd  �  EXCEPTION_ROUTINE �)�  �  �  P  �    �   PEXCEPTION_ROUTINE �   �  "_M128A j(8  	Low k�   	High l�   #M128A m  $8  Y �       2   $8  j  2   S  z  2  _ _XMM_SAVE_AREA32  ��  	ControlWord �
`   	StatusWord �
`  	TagWord �
S  	Reserved1 �
S  	ErrorOpcode �
`  	ErrorOffset �m  	ErrorSelector �
`  	Reserved2 �
`  	DataOffset �m  	DataSelector �
`  	Reserved3 �
`  	MxCsr �m  	MxCsr_Mask �m  %FloatRegisters �H   %XmmRegisters �Y  �
Reserved4 �
j  � #XMM_SAVE_AREA32 �z  &��H!  %Header �H!   %Legacy �H   %Xmm0 �8  �%Xmm1 �8  �%Xmm2 �8  �%Xmm3 �8  �%Xmm4 �8  �%Xmm5 �8  �!Xmm6 �8   !Xmm7 �8  !Xmm8 �8   !Xmm9 �8  0!Xmm10 �8  @!Xmm11 �8  P!Xmm12 �8  `!Xmm13 �8  p!Xmm14 �8  �!Xmm15 �8  � $8  Y!  2   ' ��!  (FltSave ��  (FloatSave ��  )    $8  �!  2   #CONTEXT �  PCONTEXT �  _RUNTIME_FUNCTION �%"  	BeginAddress �m   	EndAddress �m  	UnwindData �m   PRUNTIME_FUNCTION �@"  �!  ��        V"  2   EXCEPTION_RECORD �
V  PEXCEPTION_RECORD �
�"  V"  _UNWIND_HISTORY_TABLE_ENTRY �
�"    �
�   *  �
%"   UNWIND_HISTORY_TABLE_ENTRY �
�"  _UNWIND_HISTORY_TABLE ��
u#  	Count �
7   	Search �
E  	LowAddress �
�  	HighAddress �
�  	Entry �
 u#   �"  �#  2   UNWIND_HISTORY_TABLE �
�"  PUNWIND_HISTORY_TABLE �
�#  �"  DISPATCHER_CONTEXT �
&�#  _DISPATCHER_CONTEXT P�

�$  	ControlPc �
�     �
�  *  �
%"  	EstablisherFrame �
�  	TargetIp �
�   	ContextRecord �
�!  (	LanguageHandler �
�  0	HandlerData �
�  8	HistoryTable �
�#  @	ScopeIndex �
7  H	Fill0 �
7  L PDISPATCHER_CONTEXT �
'%  �#  GUID_MAX_POWER_SAVINGS �q  GUID_MIN_POWER_SAVINGS �q  GUID_TYPICAL_POWER_SAVINGS �q  NO_SUBGROUP_GUID �q  ALL_POWERSCHEMES_GUID �q  GUID_POWERSCHEME_PERSONALITY �q  GUID_ACTIVE_POWERSCHEME �q  GUID_IDLE_RESILIENCY_SUBGROUP �q  GUID_IDLE_RESILIENCY_PERIOD �q  GUID_DIS�      K_COALESCING_POWERDOWN_TIMEOUT �q  GUID_EXECUTION_REQUIRED_REQUEST_TIMEOUT �q  GUID_VIDEO_SUBGROUP �q  GUID_VIDEO_POWERDOWN_TIMEOUT �q  GUID_VIDEO_ANNOYANCE_TIMEOUT �q  GUID_VIDEO_ADAPTIVE_PERCENT_INCREASE �q  GUID_VIDEO_DIM_TIMEOUT �q  GUID_VIDEO_ADAPTIVE_POWERDOWN �q  GUID_MONITOR_POWER_ON �q  GUID_DEVICE_POWER_POLICY_VIDEO_BRIGHTNESS �q  GUID_DEVICE_POWER_POLICY_VIDEO_DIM_BRIGHTNESS �q  GUID_VIDEO_CURRENT_MONITOR_BRIGHTNESS �q  GUID_VIDEO_ADAPTIVE_DISPLAY_BRIGHTNESS �q  GUID_CONSOLE_DISPLAY_STATE �q  GUID_ALLOW_DISPLAY_REQUIRED �q  GUID_VIDEO_CONSOLE_LOCK_TIMEOUT �q  GUID_ADAPTIVE_POWER_BEHAVIOR_SUBGROUP �q  GUID_NON_ADAPTIVE_INPUT_TIMEOUT �q  GUID_DISK_SUBGROUP �q  GUID_DISK_POWERDOWN_TIMEOUT �q  GUID_DISK_IDLE_TIMEOUT �q  GUID_DISK_BURST_IGNORE_THRESHOLD �q  GUID_DISK_ADAPTIVE_POWERDOWN �q  GUID_SLEEP_SUBGROUP �q  GUID_SLEEP_IDLE_THRESHOLD �q  GUID_STANDBY_TIMEOUT �q  �      GUID_UNATTEND_SLEEP_TIMEOUT �q  GUID_HIBERNATE_TIMEOUT �q  GUID_HIBERNATE_FASTS4_POLICY �q  GUID_CRITICAL_POWER_TRANSITION �q  GUID_SYSTEM_AWAYMODE �q  GUID_ALLOW_AWAYMODE �q  GUID_ALLOW_STANDBY_STATES �q  GUID_ALLOW_RTC_WAKE �q  GUID_ALLOW_SYSTEM_REQUIRED �q  GUID_SYSTEM_BUTTON_SUBGROUP �q  GUID_POWERBUTTON_ACTION �q  GUID_SLEEPBUTTON_ACTION �q  GUID_USERINTERFACEBUTTON_ACTION �q  GUID_LIDCLOSE_ACTION �q  GUID_LIDOPEN_POWERSTATE �q  GUID_BATTERY_SUBGROUP �q  GUID_BATTERY_DISCHARGE_ACTION_0 �q  GUID_BATTERY_DISCHARGE_LEVEL_0 �q  GUID_BATTERY_DISCHARGE_FLAGS_0 �q  GUID_BATTERY_DISCHARGE_ACTION_1 �q  GUID_BATTERY_DISCHARGE_LEVEL_1 �q  GUID_BATTERY_DISCHARGE_FLAGS_1 �q  GUID_BATTERY_DISCHARGE_ACTION_2 �q  GUID_BATTERY_DISCHARGE_LEVEL_2 �q  GUID_BATTERY_DISCHARGE_FLAGS_2 �q  GUID_BATTERY_DISCHARGE_ACTION_3 �q  GUID_BATTERY_DISCHARGE_LEVEL_3 �q  GUID_BATTERY_DISCHARGE_FLAGS�      _3 �q  GUID_PROCESSOR_SETTINGS_SUBGROUP �q  GUID_PROCESSOR_THROTTLE_POLICY �q  GUID_PROCESSOR_THROTTLE_MAXIMUM �q  GUID_PROCESSOR_THROTTLE_MINIMUM �q  GUID_PROCESSOR_ALLOW_THROTTLING �q  GUID_PROCESSOR_IDLESTATE_POLICY �q  GUID_PROCESSOR_PERFSTATE_POLICY �q  GUID_PROCESSOR_PERF_INCREASE_THRESHOLD �q  GUID_PROCESSOR_PERF_DECREASE_THRESHOLD �q  GUID_PROCESSOR_PERF_INCREASE_POLICY �q  GUID_PROCESSOR_PERF_DECREASE_POLICY �q  GUID_PROCESSOR_PERF_INCREASE_TIME �q  GUID_PROCESSOR_PERF_DECREASE_TIME �q  GUID_PROCESSOR_PERF_TIME_CHECK �q  GUID_PROCESSOR_PERF_BOOST_POLICY �q  GUID_PROCESSOR_PERF_BOOST_MODE �q  GUID_PROCESSOR_IDLE_ALLOW_SCALING �q  GUID_PROCESSOR_IDLE_DISABLE �q  GUID_PROCESSOR_IDLE_STATE_MAXIMUM �q  GUID_PROCESSOR_IDLE_TIME_CHECK �q  GUID_PROCESSOR_IDLE_DEMOTE_THRESHOLD �q  GUID_PROCESSOR_IDLE_PROMOTE_THRESHOLD �q  GUID_PROCESSOR_CORE_PARKING_INCREASE_THRESHOLD �q  GUID_PROCES�      SOR_CORE_PARKING_DECREASE_THRESHOLD �q  GUID_PROCESSOR_CORE_PARKING_INCREASE_POLICY  q  GUID_PROCESSOR_CORE_PARKING_DECREASE_POLICY q  GUID_PROCESSOR_CORE_PARKING_MAX_CORES q  GUID_PROCESSOR_CORE_PARKING_MIN_CORES q  GUID_PROCESSOR_CORE_PARKING_INCREASE_TIME q  GUID_PROCESSOR_CORE_PARKING_DECREASE_TIME q  GUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_DECREASE_FACTOR q  GUID_PROCESSOR_CORE_PARKING_AFFINITY_HISTORY_THRESHOLD q  GUID_PROCESSOR_CORE_PARKING_AFFINITY_WEIGHTING q  GUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_DECREASE_FACTOR 	q  GUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_HISTORY_THRESHOLD 
q  GUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_WEIGHTING q  GUID_PROCESSOR_CORE_PARKING_OVER_UTILIZATION_THRESHOLD q  GUID_PROCESSOR_PARKING_CORE_OVERRIDE q  GUID_PROCESSOR_PARKING_PERF_STATE q  GUID_PROCESSOR_PARKING_CONCURRENCY_THRESHOLD q  GUID_PROCESSOR_PARKING_HEADROOM_THRESHOLD q  GUID_PR�      OCESSOR_PERF_HISTORY q  GUID_PROCESSOR_PERF_LATENCY_HINT q  GUID_PROCESSOR_DISTRIBUTE_UTILITY q  GUID_SYSTEM_COOLING_POLICY q  GUID_LOCK_CONSOLE_ON_WAKE q  GUID_DEVICE_IDLE_POLICY q  GUID_ACDC_POWER_SOURCE q  GUID_LIDSWITCH_STATE_CHANGE q  GUID_BATTERY_PERCENTAGE_REMAINING q  GUID_GLOBAL_USER_PRESENCE q  GUID_SESSION_DISPLAY_STATUS q  GUID_SESSION_USER_PRESENCE q  GUID_IDLE_BACKGROUND_TASK q  GUID_BACKGROUND_TASK_NOTIFICATION q  GUID_APPLAUNCH_BUTTON q  GUID_PCIEXPRESS_SETTINGS_SUBGROUP  q  GUID_PCIEXPRESS_ASPM_POLICY !q  GUID_ENABLE_SWITCH_FORCED_SHUTDOWN "q  PPM_PERFSTATE_CHANGE_GUID  q  PPM_PERFSTATE_DOMAIN_CHANGE_GUID !q  PPM_IDLESTATE_CHANGE_GUID "q  PPM_PERFSTATES_DATA_GUID #q  PPM_IDLESTATES_DATA_GUID $q  PPM_IDLE_ACCOUNTING_GUID %q  PPM_IDLE_ACCOUNTING_EX_GUID &q  PPM_THERMALCONSTRAINT_GUID 'q  PPM_PERFMON_PERFSTATE_GUID (q  PPM_THERMAL_POLICY_CH�      ANGE_GUID )q  RPC_IF_HANDLE B�  IWinTypesBase_v0_1_c_ifspec )+:  IWinTypesBase_v0_1_s_ifspec *+:  IID_IUnknown Wq  IID_AsyncIUnknown �q  IID_IClassFactory mq  IID_IMarshal nq  IID_INoMarshal Uq  IID_IAgileObject �q  IID_IAgileReference �q  IID_IMarshal2 -q  IID_IMalloc �q  IID_IStdMarshalInfo iq  IID_IExternalConnection �q  IID_IMultiQI Gq  IID_AsyncIMultiQI �q  IID_IInternalUnknown q  IID_IEnumUnknown hq  IID_IEnumString q  IID_ISequentialStream �q  IID_IStream Mq  IID_IRpcChannelBuffer �	q  IID_IRpcChannelBuffer2 ;
q  IID_IAsyncRpcChannelBuffer �
q  IID_IRpcChannelBuffer3 q  IID_IRpcSyntaxNegotiate �q  IID_IRpcProxyBuffer �q  IID_IRpcStubBuffer Vq  IID_IPSFactoryBuffer q  IID_IChannelHook �q  IID_IClientSecurity �q  IID_IServerSecurity mq  IID_IRpcOptions q  IID_IGlobalOptions �q  IID_ISurrogate !q  IID_IGlobalInterfaceTable ��      q  IID_ISynchronize q  IID_ISynchronizeHandle �q  IID_ISynchronizeEvent �q  IID_ISynchronizeContainer Aq  IID_ISynchronizeMutex �q  IID_ICancelMethodCalls q  IID_IAsyncManager �q  IID_ICallFactory q  IID_IRpcHelper fq  IID_IReleaseMarshalBuffers �q  IID_IWaitMultiple ,q  IID_IAddrTrackingControl �q  IID_IAddrExclusionControl �q  IID_IPipeByte hq  IID_IPipeLong �q  IID_IPipeDouble Jq  IID_IComThreadingInfo $q  IID_IProcessInitControl �q  IID_IFastRundown q  IID_IMarshalingStream Jq  IID_ICallbackWithNoReentrancyToApplicationSTA 	q  GUID_NULL �  CATID_MARSHALER �  IID_IRpcChannel �  IID_IRpcStub �  IID_IStubManager �  IID_IRpcProxy �  IID_IProxyManager �  IID_IPSFactory �  IID_IInternalMoniker �  IID_IDfReserved1 �  IID_IDfReserved2 �  IID_IDfReserved3 �  CLSID_StdMarshal �  CLSID_AggStdMarshal �  CLSID_StdAsyncActManager �      �  IID_IStub �  IID_IProxy �  IID_IEnumGeneric �  IID_IEnumHolder �  IID_IEnumCallback  �  IID_IOleManager !�  IID_IOlePresObj "�  IID_IDebug #�  IID_IDebugStream $�  CLSID_PSGenObject %�  CLSID_PSClientSite &�  CLSID_PSClassObject '�  CLSID_PSInPlaceActive (�  CLSID_PSInPlaceFrame )�  CLSID_PSDragDrop *�  CLSID_PSBindCtx +�  CLSID_PSEnumerators ,�  CLSID_StaticMetafile -�  CLSID_StaticDib .�  CID_CDfsVolume /�  CLSID_DCOMAccessControl 0�  CLSID_GlobalOptions 1�  CLSID_StdGlobalInterfaceTable 2�  CLSID_ComBinding 3�  CLSID_StdEvent 4�  CLSID_ManualResetEvent 5�  CLSID_SynchronizeContainer 6�  CLSID_AddrControl 7�  CLSID_CCDFormKrnl 8�  CLSID_CCDPropertyPage 9�  CLSID_CCDFormDialog :�  CLSID_CCDCommandButton ;�  CLSID_CCDComboBox <�  CLSID_CCDTextBox =�  CLSID_CCDCheckBox >�  CLSID_CCDLabel ?�  CLSID_CCDOptionButton @�  CLSID_CCDListBox A�  CLSI�      D_CCDScrollBar B�  CLSID_CCDGroupBox C�  CLSID_CCDGeneralPropertyPage D�  CLSID_CCDGenericPropertyPage E�  CLSID_CCDFontPropertyPage F�  CLSID_CCDColorPropertyPage G�  CLSID_CCDLabelPropertyPage H�  CLSID_CCDCheckBoxPropertyPage I�  CLSID_CCDTextBoxPropertyPage J�  CLSID_CCDOptionButtonPropertyPage K�  CLSID_CCDListBoxPropertyPage L�  CLSID_CCDCommandButtonPropertyPage M�  CLSID_CCDComboBoxPropertyPage N�  CLSID_CCDScrollBarPropertyPage O�  CLSID_CCDGroupBoxPropertyPage P�  CLSID_CCDXObjectPropertyPage Q�  CLSID_CStdPropertyFrame R�  CLSID_CFormPropertyPage S�  CLSID_CGridPropertyPage T�  CLSID_CWSJArticlePage U�  CLSID_CSystemPage V�  CLSID_IdentityUnmarshal W�  CLSID_InProcFreeMarshaler X�  CLSID_Picture_Metafile Y�  CLSID_Picture_EnhMetafile Z�  CLSID_Picture_Dib [�  GUID_TRISTATE \q  IWinTypes_v0_1_c_ifspec (+:  IWinTypes_v0_1_s_ifspec )+:  IID_IMallocSpy �q  IID_IBindCtx :q  �      IID_IEnumMoniker J q  IID_IRunnableObject � q  IID_IRunningObjectTable �!q  IID_IPersist i"q  IID_IPersistStream �"q  IID_IMoniker j#q  IID_IROTData X%q  IID_IEnumSTATSTG �%q  IID_IStorage X&q  IID_IPersistFile A(q  IID_IPersistStorage �(q  IID_ILockBytes �)q  IID_IEnumFORMATETC �*q  IID_IEnumSTATDATA l+q  IID_IRootStorage ,q  IID_IAdviseSink �,q  IID_AsyncIAdviseSink s-q  IID_IAdviseSink2 �.q  IID_AsyncIAdviseSink2 ./q  IID_IDataObject �/q  IID_IDataAdviseHolder 1q  IID_IMessageFilter �1q  FMTID_SummaryInformation ]2�  FMTID_DocSummaryInformation _2�  FMTID_UserDefinedProperties a2�  FMTID_DiscardableInformation c2�  FMTID_ImageSummaryInformation e2�  FMTID_AudioSummaryInformation g2�  FMTID_VideoSummaryInformation i2�  FMTID_MediaFileSummaryInformation k2�  IID_IClassActivator s2q  IID_IFillLockBytes �2q  IID_IProgressNotify �3q  IID_ILayoutStorage �3q  IID_IBloc�      kingLock �4q  IID_ITimeAndNoticeControl �4q  IID_IOplockStorage N5q  IID_IDirectWriterLock �5q  IID_IUrlMon M6q  IID_IForegroundTransfer �6q  IID_IThumbnailExtractor 7q  IID_IDummyHICONIncluder �7q  IID_IProcessLock �7q  IID_ISurrogateService H8q  IID_IInitializeSpy �8q  IID_IApartmentShutdown �9q  IID_IOleAdviseHolder �q  IID_IOleCache bq  IID_IOleCache2 )q  IID_IOleCacheControl �q  IID_IParseDisplayName <q  IID_IOleContainer �q  IID_IOleClientSite q  IID_IOleObject �q  IOLETypes_v0_0_c_ifspec �+:  IOLETypes_v0_0_s_ifspec �+:  IID_IOleWindow $q  IID_IOleLink �q  IID_IOleItemContainer �q  IID_IOleInPlaceUIWindow v	q  IID_IOleInPlaceActiveObject 
q  IID_IOleInPlaceFrame �
q  IID_IOleInPlaceObject �q  IID_IOleInPlaceSite �q  IID_IContinue �q  IID_IViewObject �q  IID_IViewObject2 *q  IID_IDropSource �q  IID_IDropTarget [q  IID_IDropSourceNotify ��      q  IID_IEnumOLEVERB vq  IID_IServiceProvider Mq  IOleAutomationTypes_v1_0_c_ifspec �+:  IOleAutomationTypes_v1_0_s_ifspec �+:  IID_ICreateTypeInfo ;q  IID_ICreateTypeInfo2 bq  IID_ICreateTypeLib �q  IID_ICreateTypeLib2 �q  IID_IDispatch �	q  IID_IEnumVARIANT �
q  IID_ITypeComp 5q  IID_ITypeInfo �q  IID_ITypeInfo2 Pq  IID_ITypeLib �q  IID_ITypeLib2 =q  IID_ITypeChangeEvents aq  IID_IErrorInfo �q  IID_ICreateErrorInfo }q  IID_ISupportErrorInfo  q  IID_ITypeFactory uq  IID_ITypeMarshal �q  IID_IRecordInfo �q  IID_IErrorLog  q  IID_IPropertyBag zq  __MIDL_itf_msxml_0000_v0_0_c_ifspec �+:  __MIDL_itf_msxml_0000_v0_0_s_ifspec �+:  LIBID_MSXML ��  IID_IXMLDOMImplementation  �  IID_IXMLDOMNode '�  IID_IXMLDOMDocumentFragment ��  IID_IXMLDOMDocument f�  IID_IXMLDOMNodeList u�  IID_IXMLDOMNamedNodeMap ��  IID_IXMLDOMCharacterData �  IID_IXMLDOMAttribu�      te ��  IID_IXMLDOMElement �  IID_IXMLDOMText ��  IID_IXMLDOMComment %�  IID_IXMLDOMProcessingInstruction ��  IID_IXMLDOMCDATASection �  IID_IXMLDOMDocumentType ��  IID_IXMLDOMNotation �  IID_IXMLDOMEntity �  IID_IXMLDOMEntityReference ��  IID_IXMLDOMParseError a	�  IID_IXTLRuntime �	�  DIID_XMLDOMDocumentEvents =
�  CLSID_DOMDocument \
�  CLSID_DOMFreeThreadedDocument `
�  IID_IXMLHttpRequest g
�  CLSID_XMLHTTPRequest �
�  IID_IXMLDSOControl �
�  CLSID_XMLDSOControl �  IID_IXMLElementCollection �  IID_IXMLDocument J�  IID_IXMLDocument2 ��  IID_IXMLElement $�  IID_IXMLElement2 ��  IID_IXMLAttribute ��  IID_IXMLError �  CLSID_XMLDocument .�  CLSID_SBS_StdURLMoniker ~�  CLSID_SBS_HttpProtocol �  CLSID_SBS_FtpProtocol ��  CLSID_SBS_GopherProtocol ��  CLSID_SBS_HttpSProtocol ��  CLSID_SBS_FileProtocol ��  CLSID_SBS_MkProtocol ��  CLSID_SBS�      _UrlMkBindCtx ��  CLSID_SBS_SoftDistExt ��  CLSID_SBS_CdlProtocol ��  CLSID_SBS_ClassInstallFilter ��  CLSID_SBS_InternetSecurityManager ��  CLSID_SBS_InternetZoneManager ��  IID_IAsyncMoniker ��  CLSID_StdURLMoniker ��  CLSID_HttpProtocol ��  CLSID_FtpProtocol ��  CLSID_GopherProtocol ��  CLSID_HttpSProtocol ��  CLSID_FileProtocol ��  CLSID_MkProtocol ��  CLSID_StdURLProtocol ��  CLSID_UrlMkBindCtx ��  CLSID_CdlProtocol ��  CLSID_ClassInstallFilter ��  IID_IAsyncBindCtx ��  IID_IPersistMoniker Pq  IID_IMonikerProp !q  IID_IBindProtocol q  IID_IBinding �q  IID_IBindStatusCallback uq  IID_IBindStatusCallbackEx �q  IID_IAuthenticate dq  IID_IAuthenticateEx �q  IID_IHttpNegotiate Aq  IID_IHttpNegotiate2 �q  IID_IHttpNegotiate3 ;	q  IID_IWinInetFileStream �	q  IID_IWindowForBindingUI 0
q  IID_ICodeInstall �
q  IID_IWinInetInfo �q  IID_IHttpS�      ecurity q  IID_IWinInetHttpInfo yq  IID_IWinInetHttpTimeouts �q  SID_BindHost 5q  IID_IBindHost ?q  IID_IInternet Mq  IID_IInternetBindInfo �q  IID_IInternetBindInfoEx &q  IID_IInternetProtocolRoot �q  IID_IInternetProtocol �q  IID_IInternetProtocolSink q  IID_IInternetProtocolSinkStackable �q  IID_IInternetSession ?q  IID_IInternetThreadSwitch Hq  IID_IInternetPriority �q  IID_IInternetProtocolInfo Nq  CLSID_InternetSecurityManager ��  CLSID_InternetZoneManager ��  IID_IInternetSecurityMgrSite �q  IID_IInternetSecurityManager iq  IID_IInternetHostSecurityManager !q  IID_IInternetZoneManager �"q  CLSID_SoftDistExt �&�  IID_ISoftDistExt �&q  IID_ICatalogFileInfo x'q  IID_IDataFilter �'q  IID_IEncodingFilterFactory �(q  GUID_CUSTOM_CONFIRMOBJECTSAFETY 3)q  IID_IWrappedProtocol A)q  IID_IGetBindHandle �)q  IID_IBindCallbackRedirect *q  IID_IPropertyStorage ��      q  IID_IPropertySetStorage q  IID_IEnumSTATPROPSTG �q  IID_IEnumSTATPROPSETSTG Dq  IID_StdOle �  GUID_DEVINTERFACE_DISK  q  GUID_DEVINTERFACE_CDROM  q  GUID_DEVINTERFACE_PARTITION  q  GUID_DEVINTERFACE_TAPE  q  GUID_DEVINTERFACE_WRITEONCEDISK  q  GUID_DEVINTERFACE_VOLUME  q  GUID_DEVINTERFACE_MEDIUMCHANGER  q  GUID_DEVINTERFACE_FLOPPY  q  GUID_DEVINTERFACE_CDCHANGER  q  GUID_DEVINTERFACE_STORAGEPORT  q  GUID_DEVINTERFACE_COMPORT  q  GUID_DEVINTERFACE_SERENUM_BUS_ENUMERATOR  q  _SCARD_IO_REQUEST !�8d  dwProtocol !�m   cbPciLength !�m   SCARD_IO_REQUEST !��c  8d  g_rgSCardT0Pci "%.Qd  g_rgSCardT1Pci "%=Qd  g_rgSCardRawPci "%LQd  IID_IPrintDialogCallback #q  IID_IPrintDialogServices #q  _Unwind_Word $02  _Unwind_Ptr $52  _Unwind_Exception_Class $=2  *�  $Bf  _URC_NO_REASON  _URC_FOREIGN_EXCEPTION_CAUGHT _URC_FATAL_PHASE2_ERROR _URC_FATAL_PHASE1_ERROR _URC_NORMAL_STOP _URC_END_OF_STACK �      _URC_HANDLER_FOUND _URC_INSTALL_CONTEXT _URC_CONTINUE_UNWIND  _Unwind_Reason_Code $L'e  _Unwind_Exception_Cleanup_Fn $WFf  Lf  \f  f  \f   bf  +_Unwind_Exception @$Z�f  exception_class $\e   exception_cleanup $] !f  private_ $`�f   �d  �f  2   _Unwind_Action $n�  _Unwind_Stop_Fn $�g  
g  f  2g  �  �f  e  \f  2g  �   8g  _Unwind_Context (E�g  cfa G�d   ra H�d  reg Ih  disp J�$    _Unwind_Trace_Fn $��g  �g  f  �g  2g  �   _Unwind_Personality_Fn $��g  �g  f  h  �  �f  e  \f  2g   �d  h  2   ,_Unwind_Backtrace �f  0�@     W      �Ei  -trace �$�g         -trace_argument ��  o   g   .  ��#  ��t.8  ��!  ��u.�  �8g  ��s/disp_context ��#  ��s0��@     �r  �h  1Rv  0 �@     �r  i  1R01w v 1w(s81w0s1w80 2-�@     *i  1R} 1Q~  3P�@     s  1Qs1Xt   4_Unwind_DeleteException ��@            ��i  -exc �4\f  �   �   5$�@     1R11Q�R  ,_Unwind_ForcedUnwind�       �f  ��@     -       �.j  -exc �1\f  9  5  -stop ��f  v  r  6�  �&�  �  �  7�@     �j  1R�R  ,_Unwind_Resume_or_Rethrow �f  ��@            ��j  -exc �6\f  �  �  0��@     <l  �j  1R�R 8��@     s  8��@     �j   9_Unwind_ForcedUnwind_Phase2 xf  `�@     U       �qk  -exc x8\f  Z  V  :stop z�f  �  �  ;�  {
�  �  �  0��@     !s  Vk  1RCCG"1Q01X11Y�  <��@     1R11QJ1w 0  4_Unwind_Resume Z�@     �       �<l  -gcc_exc Z+\f      .  \�#  ��t/ms_exc ]V"  ��s.8  ^�!  ��v0��@     �r  l  1Ru  0��@     -s  .l  1Xv 1Ys 1w u 1w(t  8��@     s   ,_Unwind_RaiseException If  ��@     A       ��l  -exc I3\f  H  B  3��@     !s  1RCCG 1Q01X11Y�   =_GCC_specific_handler ��  ��@           �co  >ms_exc �*p"  �  �  >this_frame �8�  l  b  >ms_orig_context ��!  �  �  >ms_disp �8�$  �  �  ?gcc_per �!�g  � @ms_flags �	m  �  �  @ms_code �	m  �  �  @gcc_exc �\f  r  j  A�  ��      8g  ��@gcc_action ��f  �  �  @gcc_reason �f  	  	  Bphase2 :�@     C��@     3       cn  @stop ��f  \	  Z	  D�  ��  �	  �	  <��@     1R11Q:1Yu 1w t   2N�@     �n  1R11Yu 1w t  0��@     !s  �n  1RCCG!1Q11X41Ys  2�@     �n  1R11Q11Yu 1w }  28�@     �n  1R11Q61Yu 1w }  0��@     -s  o  1Rv 1Xs 1w |  8��@     s  0��@     -s  Uo  1Rv 1Xs 1Yu 1w |  8��@     s   =_Unwind_GetTextRelBase ��d  ��@     	       ��o  ?c �12g  R =_Unwind_GetDataRelBase ��d  ��@            ��o  ?c �12g  R =_Unwind_FindEnclosingFunction ��  `�@     *       �|p  >pc �&�  �	  �	  @entry �%"  �	  �	  A  ��  �h3r�@     s  1R�R1Q�h1X0  =_Unwind_GetRegionStart ��d  P�@            ��p  ?c �12g  R =_Unwind_GetLanguageSpecificData ��  @�@     	       �	q  ?c �:2g  R E_Unwind_SetIP �0�@            �Lq  ?c �(2g  R?val �7�d  Q =_Unwind_GetIPInfo u�d   �@            ��q  ?c u,2g  R?ip_before_insn u4�  Q =_Unwin�      d_GetIP l�d  �@            ��q  ?c l(2g  R =_Unwind_GetCFA d�d   �@            �r  ?c d)2g  R E_Unwind_SetGR Z��@            ��r  >c Z(2g  6
  2
  >index Z/�  s
  o
  >val ZC�d  �
  �
  8��@     s   =_Unwind_GetGR P�d  ��@            ��r  >c P(2g  �
  �
  >index P/�  *  &  8��@     s   F�  �  %F�  �  1'F�  �  M&Gabort abort v(HL  L  %-F	  	  N P(   �  GNU C17 8.1.0 -mtune=core2 -march=nocona -g -g -g -O2 -O2 -O2 -fno-ident -fbuilding-libgcc -fno-stack-protector -fexceptions ../../../../../src/gcc-8.1.0/libgcc/emutls.c C:\mingw810\x86_64-810-posix-seh-rt_v6-rev0\build\gcc-8.1.0\x86_64-w64-mingw32\libgcc ��@     z      �  char !  long long unsigned int long long int uintptr_t K,.  wchar_t b{  short unsigned int int �  long int !  k  �  unsigned int long unsigned int unsigned char long double double float __imp___mb_cur_max s�  4  �  E  	.    _sys_errlist �&5  _sys_nerr �      �$�  
__imp___argc �  
__imp___argv �  �  �  
__imp___wargv !�  �  �  
__imp__environ '�  
__imp__wenviron ,�  
__imp__pgmptr 2�  
__imp__wpgmptr 7�  
__imp__osplatform <B  �  
__imp__osver AB  
__imp__winver FB  
__imp__winmajor KB  
__imp__winminor PB  _amblksiz 5�  __security_cookie }Y  optarg #�  optind 1�  opterr 6�  optopt :�  )    _daylight z�  _dstbias {�  _timezone |�  �  _  	.   _tzname }O  
daylight �  
timezone �  
tzname O  short int hashval_t 	*�  htab_hash 	/�  �  �  �  �   �  htab_eq 	6     �    �  �      +  +   +  htab_hash_pointer 	��  htab_eq_pointer 	��  stringop_alg �    no_stringop  libcall rep_prefix_1_byte rep_prefix_4_byte rep_prefix_8_byte loop_1_byte loop unrolled_loop vector_loop last_alg 	 e    #     
unspec_strings 
X#  
unspecv_strings 
�#  stri�      ngop_strategy ��  max ��   alg �  noalign �	�   Y  stringop_algs 4��  unknown_size �   h  ��   �  �  	.   �  processor_costs ��  add ��   lea ��  shift_var ��  shift_const ��  mult_init �&  mult_bit ��  $divide �&  (movsx ��  <movzx ��  @large_insn ��  Dmove_ratio ��  Hmovzbl_load ��  Lint_load �;  Pint_store �;  \fp_move ��  hfp_load �;  lfp_store �;  xmmx_move  �  �mmx_load P  �mmx_store P  �xmm_move �  �ymm_move �  �zmm_move �  �sse_load &  �sse_unaligned_load 	&  �sse_store 
&  �sse_unaligned_store &  �mmxsse_to_integer �  �ssemmx_to_integer �  �gather_static �  �gather_per_elt �   scatter_static �  scatter_per_elt �  l1_cache_size �  l2_cache_size �  prefetch_block �  simultaneous_prefetches �  branch_cost �  fadd �   fmul �  $f�      div �  (fabs �  ,fchs �  0fsqrt �  4sse_op "�  8addss #�  <mulss $�  @mulsd %�  Dfmass &�  Hfmasd '�  Ldivss (�  Pdivsd )�  Tsqrtss *�  Xsqrtsd +�  \reassoc_int ,�  `reassoc_fp ,�  dreassoc_vec_int ,&�  hreassoc_vec_fp ,7�  lmemcpy 3U  pmemset 3"U  xcond_taken_branch_cost 4�  �cond_not_taken_branch_cost 6�  � �  �  &  	.     �  ;  	.   +  �  P  	.   @  �  
ix86_cost :&n    
ix86_size_cost ;%  ix86_tune_indices �  ��  X86_TUNE_SCHEDULE  X86_TUNE_PARTIAL_REG_DEPENDENCY X86_TUNE_SSE_PARTIAL_REG_DEPENDENCY X86_TUNE_SSE_SPLIT_REGS X86_TUNE_PARTIAL_FLAG_REG_STALL X86_TUNE_MOVX X86_TUNE_MEMORY_MISMATCH_STALL X86_TUNE_FUSE_CMP_AND_BRANCH_32 X86_TUNE_FUSE_CMP_AND_BRANCH_64 X86_TUNE_FUSE_CMP_AND_BRANCH_SOFLAGS 	X86_TUNE_FUSE_ALU_AND_BRANCH 
X86_TUNE_ACCUMULATE_OUTGOING_ARGS X86_TUNE_PROLOGUE_USING_MOVE X86_TUNE_E�      PILOGUE_USING_MOVE X86_TUNE_USE_LEAVE X86_TUNE_PUSH_MEMORY X86_TUNE_SINGLE_PUSH X86_TUNE_DOUBLE_PUSH X86_TUNE_SINGLE_POP X86_TUNE_DOUBLE_POP X86_TUNE_PAD_SHORT_FUNCTION X86_TUNE_PAD_RETURNS X86_TUNE_FOUR_JUMP_LIMIT X86_TUNE_SOFTWARE_PREFETCHING_BENEFICIAL X86_TUNE_LCP_STALL X86_TUNE_READ_MODIFY X86_TUNE_USE_INCDEC X86_TUNE_INTEGER_DFMODE_MOVES X86_TUNE_OPT_AGU X86_TUNE_AVOID_LEA_FOR_ADDR X86_TUNE_SLOW_IMUL_IMM32_MEM X86_TUNE_SLOW_IMUL_IMM8 X86_TUNE_AVOID_MEM_OPND_FOR_CMOVE  X86_TUNE_SINGLE_STRINGOP !X86_TUNE_MISALIGNED_MOVE_STRING_PRO_EPILOGUES "X86_TUNE_USE_SAHF #X86_TUNE_USE_CLTD $X86_TUNE_USE_BT %X86_TUNE_AVOID_FALSE_DEP_FOR_BMI &X86_TUNE_ADJUST_UNROLL 'X86_TUNE_ONE_IF_CONV_INSN (X86_TUNE_USE_HIMODE_FIOP )X86_TUNE_USE_SIMODE_FIOP *X86_TUNE_USE_FFREEP +X86_TUNE_EXT_80387_CONSTANTS ,X86_TUNE_GENERAL_REGS_SSE_SPILL -X86_TUNE_SSE_UNALIGNED_LOAD_OPTIMAL .X86_TUNE_SSE_UNALIGNED_STORE_OPTIMAL /X86_TUNE_SSE_PACKED_SINGLE_INSN_OPTIMAL 0X86_TUNE_SSE_TYPE�      LESS_STORES 1X86_TUNE_SSE_LOAD0_BY_PXOR 2X86_TUNE_INTER_UNIT_MOVES_TO_VEC 3X86_TUNE_INTER_UNIT_MOVES_FROM_VEC 4X86_TUNE_INTER_UNIT_CONVERSIONS 5X86_TUNE_SPLIT_MEM_OPND_FOR_FP_CONVERTS 6X86_TUNE_USE_VECTOR_FP_CONVERTS 7X86_TUNE_USE_VECTOR_CONVERTS 8X86_TUNE_SLOW_PSHUFB 9X86_TUNE_AVOID_4BYTE_PREFIXES :X86_TUNE_USE_GATHER ;X86_TUNE_AVOID_128FMA_CHAINS <X86_TUNE_AVX256_UNALIGNED_LOAD_OPTIMAL =X86_TUNE_AVX256_UNALIGNED_STORE_OPTIMAL >X86_TUNE_AVX128_OPTIMAL ?X86_TUNE_AVX256_OPTIMAL @X86_TUNE_DOUBLE_WITH_ADD AX86_TUNE_ALWAYS_FANCY_MATH_387 BX86_TUNE_UNROLL_STRLEN CX86_TUNE_SHIFT1 DX86_TUNE_ZERO_EXTEND_WITH_AND EX86_TUNE_PROMOTE_HIMODE_IMUL FX86_TUNE_FAST_PREFIX GX86_TUNE_READ_MODIFY_WRITE HX86_TUNE_MOVE_M1_VIA_OR IX86_TUNE_NOT_UNPAIRABLE JX86_TUNE_PARTIAL_REG_STALL KX86_TUNE_PROMOTE_QIMODE LX86_TUNE_PROMOTE_HI_REGS MX86_TUNE_HIMODE_MATH NX86_TUNE_SPLIT_LONG_MOVES OX86_TUNE_USE_XCHGB PX86_TUNE_USE_MOV0 QX86_TUNE_NOT_VECTORMODE RX86_TUNE_AVOID_VECTOR_DECODE SX86_TUNE_BRANCH_�      PREDICTION_HINTS TX86_TUNE_QIMODE_MATH UX86_TUNE_PROMOTE_QI_REGS VX86_TUNE_EMIT_VZEROUPPER WX86_TUNE_LAST X �  �  	.  W 
ix86_tune_features ��  ix86_arch_indices �  "e  X86_ARCH_CMOV  X86_ARCH_CMPXCHG X86_ARCH_CMPXCHG8B X86_ARCH_XADD X86_ARCH_BSWAP X86_ARCH_LAST  �  u  	.   
ix86_arch_features ,e  
x86_prefetch_sse ;�  _dont_use_tree_here_ 
x86_mfence Y�  �  reg_class �  *�  NO_REGS  AREG DREG CREG BREG SIREG DIREG AD_REGS CLOBBERED_REGS Q_REGS 	NON_Q_REGS 
TLS_GOTBASE_REGS INDEX_REGS LEGACY_REGS GENERAL_REGS FP_TOP_REG FP_SECOND_REG FLOAT_REGS SSE_FIRST_REG NO_REX_SSE_REGS SSE_REGS EVEX_SSE_REGS BND_REGS ALL_SSE_REGS MMX_REGS FP_TOP_SSE_REGS FP_SECOND_SSE_REGS FLOAT_SSE_REGS FLOAT_INT_REGS INT_SSE_REGS FLOAT_INT_SSE_REGS MASK_EVEX_REGS MASK_REGS  MOD4_SSE_REGS !ALL_REGS "LIM_REG_CLASSES # �  �  �  	.  P �  
dbx_register_map =�  
dbx64_register_map >�  
svr4_dbx_�      register_map ?�  processor_type �  �   PROCESSOR_GENERIC  PROCESSOR_I386 PROCESSOR_I486 PROCESSOR_PENTIUM PROCESSOR_LAKEMONT PROCESSOR_PENTIUMPRO PROCESSOR_PENTIUM4 PROCESSOR_NOCONA PROCESSOR_CORE2 PROCESSOR_NEHALEM 	PROCESSOR_SANDYBRIDGE 
PROCESSOR_HASWELL PROCESSOR_BONNELL PROCESSOR_SILVERMONT PROCESSOR_KNL PROCESSOR_KNM PROCESSOR_SKYLAKE PROCESSOR_SKYLAKE_AVX512 PROCESSOR_CANNONLAKE PROCESSOR_ICELAKE_CLIENT PROCESSOR_ICELAKE_SERVER PROCESSOR_INTEL PROCESSOR_GEODE PROCESSOR_K6 PROCESSOR_ATHLON PROCESSOR_K8 PROCESSOR_AMDFAM10 PROCESSOR_BDVER1 PROCESSOR_BDVER2 PROCESSOR_BDVER3 PROCESSOR_BDVER4 PROCESSOR_BTVER1 PROCESSOR_BTVER2  PROCESSOR_ZNVER1 !PROCESSOR_max " 
ix86_tune 	K  
ix86_arch 	K  
ix86_preferred_stack_boundary 		�  
ix86_incoming_stack_boundary 
	�  �  �  	.  P �  
regclass_map 	�  pthread_once_t ��  pthread_key_t ��  pthread_mutex_t +  
_pthread_key_dest #    __gthrea�      d_key_t 0�  __gthread_once_t 1�  __gthread_mutex_t 2�  word !.  pointer ".  (�  offset )}  ptr *+   __emutls_object  $  h  &p   align 'p  loc +�  templ ,	+   __emutls_array /8  h  1}   data 2
8   -  G  .   emutls_mutex <V  	��L     emutls_key >%  	��L     emutls_size ?}  	x�L      __emutls_register_common ���@     *       �   !obj �3   R"h  �p  Q!align �p  X!templ �#+  Y �  #__emutls_get_address +  �@     �      ��#  $obj /   m  c  %offset �}  �  �  %arr ��#  �  n  %ret �	+  X  P  &`   �!  once �=  	p�L     ''  c�@     �   �!  (3'  �  �  (#'  �  �  )v�@     g'  *R	p�L     *Q	��@       '�%  v�@     �   �[!  (&      )��@     t'  *R	��L       +�%  ��@        �(�%  @  >  )��@     �'  *R	��L        &P  *"  ,h  �}  n  l  'F&  ��@     �  ��!  (y&  �  �  (j&  �  �  )��@     �'  *Qs   -��@     �'  "  *Rt!*Q8 .��@     ��      '   /0�@     U       #  %orig_size �}  �  �  ,h  �}      0F&  r�@     r�@            ��"  (y&  �  �  (j&  �  �  )��@     �'  *Qs   -P�@     �'  �"  *Rs *Q| 3$# )r�@     �'  *R	v 3$s "#*Q0*X| 3$  '�&  &�@     0   � @#  (�&  �  �  .1�@     �'   +�#  ��@     �  �($      1�  2$  a  [  2$  �  �  -��@     �'  �#  *Rt v "# -�@     (  �#  *Xv  -��@     �'  �#  *Rv )��@     �'  *Q0      3emutls_alloc ]+  )$  4obj ]'   5ptr _	+  5ret `	+   6emutls_init R��@     4       �%  '&  ��@         U�$  (8&  �  �  )��@     *(  *R	��L     *Q0  0�&  ��@     ��@            W�$  (�&  )  '  (�&  W  U  )��@     7(  *R	��L     *Q	��@       .�@     �'   6emutls_destroy B��@     ?       ��%  $ptr B+  �  �  %arr D�#  �  �  ,h  E}  S  Q  %i F}  z  v  .��@     D(  7��@     D(  *R�R  8__gthread_mutex_unlock �  �%  9�  ,�%   V  8__gthread_mutex_lock ��  &  9�  �*�%   :__gthread_mut�      ex_init_function �F&  9�  �3�%   8__gthread_setspecific ��  �&  ;__key �(%  ;__ptr �;�   8__gthread_getspecific �+  �&  ;__key �(%   8__gthread_key_create ��   '  ;__key �( '  ;__dtor �6   %  8__gthread_once ��  D'  ;__once �#D'  ;__func �2.   =  <__gthread_active_p +�  =[  [  *=m  m  S=�  �  U=�  �  '>calloc calloc �>abort abort v(>realloc realloc �?memset __builtin_memset  =�  �  &>malloc malloc �?memcpy __builtin_memcpy  =�  �  W=�  �  $>free free �                                                                                                                                                                                           %   I  $ >  & I   :;9I   :;9I   I  :;9  	:;9  
 :;9I8   :;9I8   :;9I8   <  :;9  I  ! I/  :;9   :;9I8  9:;  9�      :;9�  :;9  :;9   I8  .?:;9n<d   I4   I   :;9I2  :;9   :;9I   :;9I?2<   I8   .?:;9n<d  !.?:;9nI<d  ".?:;9nI<d  #.?:;9n<d  $.?:;9nI<d  %.?:;9nI<d  &.?:;9n<  '.?:;9n<  (.?:;9nI<  ).?:;9n2<d  *.?:;9n2<cd  +.?:;9n2<d  ,.?:;9nI2<d  -.?:;9nI2<d  . :;9I2  // I  0/ I  1: :;9  2 :;9  3 :;9  4.?:;9n<c�d  54 :;9nI?<  69:;9  7:;9  8.?:;9n<cd  9.?:;9n2<d  :.?:;9nI2<d  ;.?:;9n2<d  <.?:;9nI2<cd  =.?:;9nI2<d  >.?:;9n�<  ? <  @ :;9I?<l  A :;9I  B/ I  C0 I  D9 :;9  E>I:;9  F(   G4 :;9I<
l  H9 :;9  I :;9I  J.?:;�      9nI<  K. ?:;9nI<  L I82  M.?:;9n2<d  N.?:;9nI2<d  O9 :;9�  P: :;9  Q<  R:;92  S :;9I?<  T4 :;9I<  U.?:;9nI<  V:;9  W9:;9  X9 :;9�  Y :;9I?<  Z.?:;9n<  [. ?:;9nI<  \:;9  ] :;9I82  ^ :;9I2  _4 :;9I?<  `.?:;9I<  a.:;9I<  b   c. ?:;9I<  d.:;9I<  e.?:;9I<  f   g I  h;   iB I  j4 G  k. ?:;9I<  l!   m   n  o4 :;9I?<  p&   q:;9n  rI  s.?:;9<  t4 G  u4 nG  v4 nG  w4 nG  x4 nG  y4 nG  z. 4@�B  {.4@�B  | :;9I  }. ?:;9I@�B   %   I  $ >  & I   :;9I   :;9I   I  :;9  	:;9  
 :;9I8   :;9I8   :;9I8   <  :;9  I  ! I/  :;9  �       :;9I8  9:;  9:;9�  :;9  :;9   I8  .?:;9n<d   I4   I   :;9I2  :;9   :;9I   :;9I?2<   I8   .?:;9n<d  !.?:;9nI<d  ".?:;9nI<d  #.?:;9n<d  $.?:;9nI<d  %.?:;9nI<d  &.?:;9n<  '.?:;9n<  (.?:;9nI<  ).?:;9n2<d  *.?:;9n2<cd  +.?:;9n2<d  ,.?:;9nI2<d  -.?:;9nI2<d  . :;9I2  // I  0/ I  1: :;9  2 :;9  3 :;9  4.?:;9n<c�d  54 :;9nI?<  69:;9  7:;9  8.?:;9n<cd  9.?:;9n2<d  :.?:;9nI2<d  ;.?:;9n2<d  <.?:;9nI2<cd  =.?:;9nI2<d  >.?:;9n�<  ? <  @ :;9I?<l  A :;9I  B/ I  C0 I  D9 :;9  E>I:;9  F(   G4 :;9I<
l  H9 :�      ;9  I :;9I  J.?:;9nI<  K. ?:;9nI<  L I82  M.?:;9n2<d  N.?:;9nI2<d  O9 :;9�  P: :;9  Q<  R:;92  S :;9I?<  T4 :;9I<  U.?:;9nI<  V:;9  W9:;9  X9 :;9�  Y :;9I?<  Z.?:;9n<  [. ?:;9nI<  \:;9  ] :;9I82  ^ :;9I2  _4 :;9I?<  `.?:;9I<  a.:;9I<  b   c. ?:;9I<  d.:;9I<  e.?:;9I<  f   g I  h;   iB I  j4 G  k. ?:;9I<  l!   m   n  o4 :;9I?<  p&   q:;9n  rI  s.?:;9<  t4 G  u4 nG  v4 nG  w4 nG  x4 nG  y4 nG  z. 4@�B  {.4@�B  | :;9I    %   %  $ >  & I   :;9I   I  4 :;9I?<   '  I  	! I/  
4 :;9I?<  'I   I  &   >I:;9  (   !   :;9   :;9�      I8  :;9   :;9I8   :;9I8  >I:;9   <  4 G:;9   %  $ >  & I   :;9I   :;9I   I  :;9   :;9I8  	 :;9I8  
 :;9I8   <  :;9  :;9  I  ! I/  4 :;9I?<  4 :;9I?<  '   I  'I  &      >I:;9  (   !   :;9   :;9I8  :;9   <  >I:;9  �:;9    I�8  ! :;9I�8  "�:;9  # :;9I�  $I�  % :;9I�8  &�:;9  '�:;9  ( :;9I�  ) I�  *>I:;9  +�:;9  ,.?:;9'I@�B  - :;9I�B  .4 :;9I  /4 :;9I  0��1  1�� �B  2��  3��1  4.?:;9'@�B  5���B  6 :;9I�B  7���B1  8�� 1  9.:;9'I@�B  :4 :;9I�B  ;4 :;9I�B  <�� �       =.?:;9'I@�B  > :;9I�B  ? :;9I  @4 :;9I�B  A4 :;9I  B
 :;9  C  D4 :;9I�B  E.?:;9'@�B  F. ?<n:;9  G. ?<n:;9  H. ?<n:;9   %  $ >  & I   :;9I   I  4 :;9I?<   '  I  	! I/  
4 :;9I?<  'I   I  &   '     >I:;9  (   !   :;9   :;9I8   :;9I8  :;9   :;9I8   :;9I8  >I:;9   <   :;9I  :;9   :;9I  ! I  4 :;9I   .?:;9'@�B  ! :;9I  " :;9I  #.?:;9'I@�B  $ :;9I�B  %4 :;9I�B  &U  '1R�BUXYW  ( 1�B  )��1  *�� �B  +1R�BUXYW  ,4 :;9I�B  -��1  .�� 1  /  01R�BXYW  1U  24 1�B  3.:;9'I   4 :;9I  54 :;9I  6.:;9'�      @�B  7���B1  8.:;9'I   9 :;9I  :.:;9'   ; :;9I  <. :;9'I   =. ?<n:;9  >. ?<n:;9  ?. ?<n:;                                                                                                                                  �  �      F:/debug/ClionWork/EFS/OS D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++ D:/MinGW-w64/mingw64/x86_64-w64-mingw32/include D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/bits D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/x86_64-w64-mingw32/bits D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/debug D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/ext F:/debug/ClionWork/EFS  main.cpp   iostream   crtdefs.h   locale.h   basic_string.h   stringfwd.h   cwchar   new   exception_ptr.h   c++config.h   type_traits   cpp_type_traits.h   stl_pair.h   debug.h   char_traits.h   cstdint   cloc�      ale   allocator.h   cstdlib   cstdio   alloc_traits.h   initializer_list   system_error   ios_base.h   cwctype   iosfwd   std_abs.h   stl_iterator_base_types.h   predefined_ops.h   new_allocator.h   numeric_traits.h   alloc_traits.h   stl_iterator.h   wchar.h   swprintf.inl   string.h   stdint.h   stdio.h   ctype.h   process.h   pthread.h   atomic_word.h   stdlib.h   malloc.h   io.h   wctype.h   excpt.h   minwindef.h   guiddef.h   winnt.h   rpcdce.h   stdlib.h   wtypesbase.h   unknwnbase.h   objidlbase.h   cguid.h   wtypes.h   objidl.h   oleidl.h   servprov.h   oaidl.h   msxml.h   urlmon.h   propidl.h   oleauto.h   winioctl.h   winsmcrd.h   winscard.h   commdlg.h   utilities.h   <built-in>      	P@     �Y.�YY� f��.� f� ��tt� �   �  �      D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++ F:/debug/ClionWork/EFS/OS/VHD D:/MinGW-w64/mingw64/x86_64-w64-mingw32/include D:/MinGW-�      w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/bits D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/x86_64-w64-mingw32/bits D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/debug D:/MinGW-w64/mingw64/lib/gcc/x86_64-w64-mingw32/8.1.0/include/c++/ext F:/debug/ClionWork/EFS  iostream   disk.h   crtdefs.h   locale.h   basic_string.h   stringfwd.h   cwchar   new   exception_ptr.h   c++config.h   type_traits   cpp_type_traits.h   stl_pair.h   debug.h   char_traits.h   cstdint   clocale   allocator.h   cstdlib   cstdio   alloc_traits.h   initializer_list   system_error   ios_base.h   cwctype   iosfwd   std_abs.h   stl_iterator_base_types.h   predefined_ops.h   new_allocator.h   numeric_traits.h   alloc_traits.h   stl_iterator.h   wchar.h   swprintf.inl   string.h   stdint.h   stdio.h   ctype.h   process.h   pthread.h   atomic_word.h   stdlib.h   malloc.h   io.h   wctype.h   excpt.h   minwindef.h   guiddef.h   winnt.�      h   rpcdce.h   stdlib.h   wtypesbase.h   unknwnbase.h   objidlbase.h   cguid.h   wtypes.h   objidl.h   oleidl.h   servprov.h   oaidl.h   msxml.h   urlmon.h   propidl.h   oleauto.h   winioctl.h   winsmcrd.h   winscard.h   commdlg.h   utilities.h   <built-in>      	@     � �G.� f9�Gtt� w    O   �      ../../../../../src/gcc-8.1.0/libgcc/config/i386  cygwin.S     	 �@     � ""gY0uKgg0=L"" �   �  �      C:/mingw810/x86_64-810-posix-seh-rt_v6-rev0/mingw64/mingw/include C:/mingw810/src/gcc-8.1.0/include ../.././gcc C:/mingw810/src/gcc-8.1.0/gcc/config/i386 C:/mingw810/src/gcc-8.1.0/libgcc ../../../../../src/gcc-8.1.0/libgcc  crtdefs.h   stdlib.h   malloc.h   process.h   getopt.h   time.h   hashtab.h   insn-constants.h   i386.h   i386-opts.h   libgcc2.h   gbl-ctors.h   libgcc2.c    T   �  �      ../../../../../src/gcc-8.1.0/libgcc C:/mingw810/x86_64-810-posix-seh-rt_v6-rev0/mingw64/mingw/include C:�      /mingw810/src/gcc-8.1.0/include ../.././gcc C:/mingw810/src/gcc-8.1.0/gcc/config/i386  unwind-seh.c   crtdefs.h   stdlib.h   malloc.h   process.h   getopt.h   time.h   hashtab.h   insn-constants.h   i386.h   i386-opts.h   excpt.h   winnt.h   minwindef.h   ctype.h   basetsd.h   guiddef.h   rpcdce.h   wtypesbase.h   unknwnbase.h   objidlbase.h   cguid.h   wtypes.h   objidl.h   oleidl.h   servprov.h   oaidl.h   msxml.h   urlmon.h   propidl.h   oleauto.h   winioctl.h   winsmcrd.h   winscard.h   commdlg.h   ./unwind.h    errhandlingapi.h     	`�@     �K~\�kYJ�?�}JKZ<YVf 	��@     KZ<YVf 	 �@     =�K�Igl	K��� J/fK2K�=! X0 . Y=W/�����	=v.
�	xf0J�+PdT���Yf�      �X�Z?
[
�$WK$8K$�H�
 � � � < .�f#JJu.JXX<X�?7]X)�X�
[
]�[*VK	&wf	XxXIK$MzJu$K$Kt��XJtX<<�� JY1b\T=XJ?+?���oAXt��g"�yX@z]��Z"O"�Y"�"�h�tKu[WX	f�KL
X 	�@     
JY�=�/z�BY�Vz<C�=��<eX�~���Y#��"t��G�UzzfP
<N
�k�#=,JfMX
J	YX.	zf �   �  �      ../../../../../src/gcc-8.1.0/libgcc C:/mingw810/x86_64-810-posix-seh-rt_v6-rev0/mingw64/mingw/include C:/mingw810/src/gcc-8.1.0/include ../.././gcc C:/mingw810/src/gcc-8.1.0/gcc/config/i386  emutls.c   ./gthr-default.h    crtdefs.h   stdlib.h   malloc.h�         process.h   getopt.h   time.h   hashtab.h   insn-constants.h   i386.h   i386-opts.h   pthread.h   <built-in>      	��@     � u=7A
.0
XY � J^=fX 	��@     L��|���z�
.�{LW( ���~Ls<<.�
��{
�<<�{	.*<�	J=��SJ��|��X�{��|���{K
���|��{�K
;=
h
��{f=�
�X�{�
J<
��
�FY	<=M
K;��@=>m�Y;Ju
�;=
0=Y;��
�X�{�
Z=Jf+�u�c��( �Z=�gK XZK                                                    �                                                                                                                                                                                                                                                                                                                                                                         ���� x �      $       P@     ?       A�Cz�   $       �@            A�CV�   $       �@     <       A�Cw�   $       �@            A�CY�      ���� x �      $   �   @            A�CV�   $   �   +@     <       A�Cw�   $   �   g@            A�CY�      ���� x �      ,   H   �@     2       A�A�n�A�         ���� x �         �  `�@     U       D@P $   �  ��@            D0Q
A       $   �  ��@            D0Q
A          �   �@               �  �@               �   �@               �  0�@               �  @�@     	          �  �      P�@            $   �  `�@     *       D@^
AF       �  ��@               �  ��@     	       \   �  ��@           B�B�A �A(�A0�A8�D��
8A�0A�(A� A�B�B�D       $   �  ��@     A       A�D0zA� ,   �  �@     �       A�A�A �A(�G�   �  ��@            D0        �  ��@     -          �  �@            l   �  0�@     W      B�B�B �B(�A0�A8�A@�AH�	G�+
HA�@A�8A�0A�(B� B�B�B�F       ���� x �      <   x  ��@     ?       A�A�A �D@p A�A�A�       $   x  ��@     4       D0i
A       L   x  �@     �      B�A�A �A(�A0�DPB
0A�(A� A�A�B�A    x  ��@     *                                                                                                                                                                       size_type vswprintf replace const_iterator __value allocator _M_local_data _Value compare _Iterator _M_get_allocator nothrow_t operator-- find_l�      ast_not_of refcount operator-= operator-> basic_string append piecewise_construct_t iterator __is_signed _Traits _M_current __max_digits10 find_last_of deallocate operator* operator+ operator- char_type length to_char_type operator= new_allocator find_first_of rfind to_int_type allocate __normal_iterator const_pointer operator++ operator[] _CharT insert value_type assign operator+= find _S_copy_chars __max _Alloc_hider _Container reference __digits10 const_reference int_type swprintf __min eq_int_type exception_ptr difference_type find_first_not_of pointer max_size initializer_list _Alloc __max_exponent10 __digits allocator_type size_type vswprintf replace const_iterator __value allocator _M_local_data _Value compare _Iterator _M_get_allocator nothrow_t operator-- find_last_not_of refcount operator-= operator-> basic_string append piecewise_construct_t iterator __is_signed _Traits _M_current __max_digits10 find_last_of deallocate operator* operator+ operator- char_type length to_char_type operator= ne�      w_allocator find_first_of rfind to_int_type allocate __normal_iterator const_pointer operator++ operator[] _CharT insert value_type assign operator+= find _S_copy_chars __max _Alloc_hider _Container reference __digits10 const_reference int_type swprintf __min eq_int_type exception_ptr difference_type find_first_not_of pointer max_size initializer_list _Alloc __max_exponent10 __digits allocator_type ../../../../../src/gcc-8.1.0/libgcc/config/i386/cygwin.S C:\mingw810\x86_64-810-posix-seh-rt_v6-rev0\build\gcc-8.1.0\x86_64-w64-mingw32\libgcc GNU AS 2.30 RtlLookupFunctionEntry stop_argument gcc_context RtlCaptureContext RtlVirtualUnwind RtlUnwindEx ImageBase ms_history FunctionEntry ms_context refcount RaiseException pthread_once size pthread_mutex_lock pthread_getspecific pthread_key_create pthread_setspecific __mutex pthread_mutex_init pthread_mutex_unlock                              �      �       R�             _             �R�      '       _                        �      [      �       Q[             ^             �Q�      '       ^                        �      �       R�      �       Q�      �       �R��      �       R                    �      �       R�      �       �R�                    �      �       Q�      �       �Q�                    �      �       X�      �       �X�                        `      o       Ro      u       �R�u      y       Ry      |       �R�                                    R                y                   &       ;        p                     &       ;        p0;       H        QH       J        �h                    �      �       R�      _       S                      `             R      �       Q�      �       y                                   P      �       R�      1       S1      ;       R;      E       SE      M       �R�M      a       Ra      *       S*      @       R@      Q       S                          P      u  �           Qu      H       VH      M       �Q�M      X       QX      Q       V                                  P      �       X�      1       \1      ;       X;      J       \J      M       �X�M      �       X�      *       \*      =       X=      Q       \                                      P      �       Y�      1       �Y�1      ;       T;      M       �Y�M      j       Tj      r       Yr      �       ���      �       �Y��      %       T%      *       �Y�*      Q       T                                  _      �       P1      ;       PM      T       PT      a       ra      e       Pe      w       s�      �       P*      .       P.      :       r                                   _      �       r �      �       Q1      ;       QM      a       r a      o       Qo      w       s �      �       Q�      �       s *      5       Q5      :       r                      �        _      �       r �      ;       UM      a       r a      Q       U                   �      �       Qa      �       :�                      �             P�      �       P�      �       P                 a      w       u                   a      w       u0w      �       P                                  R      *       �R�                                 P#      %       P                    �       �        R�       �        �R�                    �       �        Q�       �        �Q�                    �       �        X�       �        �X�                    `       {        R{       |        �R�                    `       {        Q{       |        �Q�                          �       �        R�       �        U�       �        �R��       �        R�       H       U                            �       �        T�       H       T�      �       T             T      "       u"      +       T          �                                �       �        P�       �        S             P      (       S(      >       P>      D       S�      �       P�      �       S�      �       P�      �       S                       �       �        YD      ^       Y�      �       Y�      �       Y                 �       �       
 ��@     �                 �       �       
 p�L     �                 �       �       
 ��L     �                 �             
 ��L     �                  "      D       V                   7      >       P>      D       S                 7      >       R                 �      �       V                      �      �       \�      �       p �      �      ) t v 1$t #���������v 1$#���������+( �                 �      �       S                 �      �      	 ��L                      �       �       	 ��L                         D      �       U�             U+      B       U                     �       _      �       P�             P+      9       P                      s      �       Y
             Y+      9       Y                 D       R       
 ��L     �                 R       e       
 ��@     �                 R       e       
 ��L     �                                        R       9        T9       >        R>       ?        �R�                                      R       9        T9       >        R>       ?        �R�                  
       :        U                   
               0�       0        S                                                                                                                                                                                                                                                                                                                                                               D       D       D       R                       �       �       �       �               �              �       �       �       �       �       �       �                   0                      �       �       �       �                       �       �       �       �                       �       �       �                                   D      B      H                      .      4      7      D                      D      �      �            0      B                                      .file   M   ��  gcrtexe.c              j                                �              �   �U                        �   �U                        �   �U                          �U                        )  @T                        G  pU                        e             p  0U                        �  �H                        �  0          �  `U                    envp           argv           argc                �              �   U                        �  �            �T     �                         3  �T                        Y             c   T                        �  �T                        �  PT                    mainret            �  �T                        �  �T                        �  U                           U                        )  �          ;  �      .l_endw �          E  �      .l_start�      .l_end  �      atexit            T  @U                        z  PU                    .text          )  K             .data                           .bss           $                 .xdata         p   
             .pdata         T                    �                            �                         .file   \   ��  gcygming-crtbegin.c    �  0                           �  @      .text   0                     .data                           .bss    0                        .xdata  p           �                  .pdata  T                      .file   �   ��  gmain.cpp              �              �  0       main    P                           �  �N                          �N                    __tcf_0 �          _  �          �  �      .text   P     �                .data                           .bss    0                       .rdata                          .xdata  x      0                 .pdata  l      0                .ctors  (�	                        �         c�  &                �                             �      
   0                    �                            �                             �  ��     ?                     �         �                .file   �   ��  gdisk.cpp              �             �  @       __tcf_0                            _  +          �  g      .text        u                .data                           .bss    @    �                         .rdata                         .xdata  �      $                 .pdata  �      $   	             .ctors  0�	                        �  c�     L�  %                �       �                    �  0   
   0                    �       �                   �                           �  ��     ?                     �  �      �                .text   �      .data          .bss    P       .idata$7       .idata$5d      .idata$4�      .idata$6�      .text   �      .data          .bss    P       .idata$7�      .idata$5�      .idata$4�      .idata$6�      .text   �      .data          .bss    P       .idata$7�      .idata$5�      .idata$4�      .idata$6t      .text   �      .data          .bss    P       .idata$7|      .idata$5      .idata$4�       .idata$6D
      .file   �   ��  gfake              hname   <       fthunk  �      .text   �         �                    .data                           .bss    P                        .idata$2                       .idata$4<       .idata$5�      .file   Kj  ��  gfake              .text   �                       .data                           .bss    P                        .idata$4�                      .idata$5l                      .idata$7$                      .text   �                       .data                           .bss    P                                    �                     8  `     �                     \  �     �                     �  `     P                     �        P                     �  �     P                       �     �                     %        �                     H  �     �                     l  @     P                     �  �     P                     �  �     P                     �  �+                         �  �*               �                   -                           �)                         ,  `'                         <  @&                         L  �(                         \   %                         k  0P	                          �  pM                        �  �M                        �  0I                        !  PQ                        ]   O                        �  I                        �   I                        	  P                        !	  `N                        9	   P                        O	  pN                        h	  �N                        �	  `I                        �	  `Q                        �	  O                        :
  @I                        m
  PI                        �
  �N                        �
   Q                        �
  �N                          �P                      �        H  �N                        b  �N                        |  �S                        �  �S                        �  0P	         �  �W	           �W	         .  �L	         P  �I                        }  pI                        �  �I                        �  �I                          �I                        1  �I                    .text   �                       .data                           .bss    P                            _  0P	    �  M                 }  �                          �  �                          �  �W	    �                    �  L                          �  �                            �L	    g  8                 ?  l     )                    h  �                          �  ��                       �  ��                          �  ��                       /  ��         a  ��         x  ���               �  ��         �  `�     __tcf_0 ��	         �  `.            ��                       C  ��         o  0�     (                   �  ��    $                   �  ��         �  p�                       3  p�         a  ��     (                   �  @�    $                   �  @�         �  �    S                     �         ?  �d                        s  �         �  �         �   �         �   �         �  pZ         �  �K                          �r         .  ��         T  �U          ^  �         �  Ч         �  ��         �  ��         �  �         �  �         �  �           `�         (  `�         D  @Z         ]  ��         �  �K                        �  Г         �   �         5  ��         h  p          �  @d                        �  ��                                �  �                          ��                         +  �l                        H  ��     '                    z   �     )                    �  �                     .text   �                       .data                           .bss    P                        .rdata         �                     �  �                           �                         9  �                         r  �                         �  ��                         �  �                          �  �                            ��                        !  �                          ?                           ]  `�                        �  �                          �                           �  ��	                        �  �                          	                              �                         K  ,                        ~        �                         �  8                        �  �                           D                        N  �                         �  P                        �  �                        �  \                          �                         "  �                          =  h                         X   �                         y  �                          �  t                         �  pZ    5                   �  �     ,                      �                         %  �r    (  	                 @       -                    \  �                         x  ��    A                    �  L                          �  �                         �  �    #                    *  T                          W  �                         �  Ч                        �  \                          �  �                                 ��    1  
                 !  `     =                    ?  �                         ]  �    T                    w  �                          �  �                         �  �    )                    �  �                          �  �                         �  `�    �                     �     0                    9  �                         \  @Z    *                    {  �                          �  �                         �  ��    .                   �  �     �                    >   �                         �   Г    H                    �   h                          �                            0!   �    ?                    o!  p                          �!                           �!  ��    �  !                 ("  |     9                    b"                           �"  �U                                �"  P"                          �"  p"                          �"  0[                          #  `"                          ?#  �"                          [#  �"                          y#  @"                          �#  @Y                          �#  `[                          �#  p[                          �#  `Y                          $  @[                          %$  P[                          B$   [                          ]$  PY                          w$  p                          �$  `.                          �                                /           __tcf_0 ��	         	%  0.          C               3               �               �               ?%  ��         e%  P          �%  ��    /                   �%  ��                        &   �         &  �          7&  �          T&  �          p&             �&  @          �&  PK                              �&  @          �&  �L                        
'  �Q                        5'  `          Z'             y'  �O                        �'  @L                        �'  �R                        (  P          <(   M                        �(  �R                        �(  p          �(  @M                        F)  `O                        q)  �          �)   L                        �)  �Q                        �)             *  �          5*   O                        h*  �K                        �*   R                        �*  �          �*  �          +  0O                        J+  �K                        ~+  �O                        �+  �          �+  �L                        Q,  �O                        �,  �          �,  �L                        $-  �Q                        P-  �                v-  �          �-  `J                        �-  �O                        .  @          6.  `L                        �.  PS                        �.  `          �.  �M                        M/  �          l/   L                        �/  �          �/  `K                        �/  `          �/  �L                        0  �Q                        D0             i0             �0  �O                        �0  PL                        �0  �R                        .1  `          K1  0M                        �1  �R                        �1  �          2  PM                        U2  pO                        �2  �          �2  L                        �2  R                        �2             "3             D3  @O                        w3  �K                        �3   R                        �3  �          4                   &4  PO                        Y4  �K                        �4  �O                        �4  �          5  �L                        `5  �O                        �5  �          �5  �L                        36  �Q                        _6  �
          �6             �6  pJ                        �6  �O                        &7  P          E7  pL                        �7  `S                        �7  p          8   N                        \8  �          {8  0L                        �8  �R                        �8  �          �8  �L                        9  �R                        79  �          W9  �L                        ~9   �         �9  P�         �9  �          �9  pK                        :  �K                        *:  ��         H:  �K                        m:   �         ~:   �         �:  Щ               �:  `          �:  ��     .text   �                       .data                           .bss    P                        .rdata  �      P                     �  ��	                        �  �                         	  (                         �:  ��    {                    ;  �                         4;  4                         a;  �                         �;  @                        �;   �    �  �                �;  �     �                    
<  L                         (<  P�    5                    Q<  |                          {<  X                         �<  ��    [                    �<  �                          �<  d                         =   �    �                    *=  �     -                    B=  p                         Z=  Щ    +                    w=  �                          �=  |                         �=  ��                             �=  �     =                    �=  �                         >   X                         :>  �Z     8                    j>  `Z                         �>  �Z     H                    �>  �Y     8                    �>   Z                         ?   Z     8                    ;?  �Y     8                    c?  �
     �                    �?        �                     �?  �     �                     �?        �                     @  �     �                    B@        p                     p@  �     p                     �@  `     �                     �@  �                          �@  �                          A  �                           :A  p                          _A  P                          �A        (                     �A  �                          �A  �                          �A                             B        	                           FB  `                          iB  �                          �B  `                          �B                             �B  �                          �B  �     �                    C  �                           =C  `                          bC  @                          �C  �     (                     �C  �                          �C  �                          �C  �                          !D  �                          ID  @                          lD  p                          �D  P                          �D                             �D  �                          �D  @     @                    E  �     p                    >E  �     p                    aE                             �E  �     0                     �E  `                          �E  �     (                     �E  P                          +F  0.            
                    gF  0�                          �F   J                        �F  J                        	G  p�         JG  ��         oG  ��         �G  p�         �G  �         �G  �         H  ��         (H  ��         iH  �         �H  @�         �H  @�         �H  �         I  p�         >I  p�         cI  @�     .text   �                       .data                           .bss    P                        .rdata  0                          �I  0�    U                   �I                            J  �                         _J  p�    U                   �J                            �J  �                         6K  ��    H                    aK                            �K  �                         �K  p�    0                    �K  4                         L  �                         <L  �    H                    gL  P                                �L  �                         �L  ��    0                    �L  p                         M  �                         BM  ��    f                   �M  �                          �M  �                         N  �    f                   `N  �                          �N  �                         �N  @�    H                    O  �                          GO  �                         sO  �    0                    �O  �                         �O                            �O  p�    H                    !P  �                          MP                           yP  @�    0                    �P  �                         �P                           �P  �h    ]                   'Q  �h                          LQ  ��                         uQ  ph    0                   �Q  ph         �Q  �a    ]                   �Q        �a         R  ��                         >R  �a    0                   iR  �a         �R  @w    ]                   �R  @w         �R  0�                         S  w    0                   2S  w         WS  �o    ]                   �S  �o         �S  �                         �S  �o    0                   �S  �o          T  ��         LT  p�         �T  ��         �T  ��         �T  @P                        U  ��         !U  ��         >U   �         [U  0P                        �U   �         �U  ��         �U   �         �U  0�         0V  ��         MV  `P                        vV  ��         �V  P�         �V  ��         �V  PP                        �V  ��         W  ��         0W  ��                         YW  z                        �W  ��                         �W  �y                        �W  ��                               �W  Pz                        &X  ��                         OX  0z                    .text   �                       .data                           .bss    P                            xX                           �X  $                        �X                          �X  0                        (Y  8                         TY  <                        �Y  @                        �Y  H                        �Y  \                         Z  T                        0Z  d                        \Z  `                        �Z  �                         �Z  l                        �Z  �                        [  x                        8[  ��    
                    j[  �                          �[  �                     .rdata  @                          �[  p�    Q                   \  �                                O\  �                         �\  ��    Q                   �\  �                          ]  �                         N]  ��    H                    q]  �                          �]  �                         �]  ��    0                    �]  �                          ^  �                         $^   �    H                    G^  �                          k^  �                         �^  ��    0                    �^                           �^  �                         �^   �    b                   9_  0                          y_  �                         �_  0�    b                   �_  8                          8`  �                         x`  ��    H                    �`  @                          �`  �                         �`  P�    0                    a  `                         *a  �                         Na  ��          H                    qa  |                          �a                           �a  ��    0                    �a  �                          b                           $b  @8	                          Yb  �I                        �b  �I                        �b  �;	         �b  �;	         �b  P;	         c  �;	         Gc  �>	         ec  �>	         �c  �>	     .text   �                       .data                           .bss    P                        .rdata  P     "                     �c  @8	    /                   �c  �                          d                            Td  �;	    H                    xd  �                          �d  ,                         �d  P;	    0                    �d  �                         e  8                         0e  �;	                       ke  �                          �e  D                               �e  �>	    H                    f                            ,f  P                         Qf  �>	    0                    uf  $                         �f  \                         �f  �<    R                   �f  �<                          g  `�                         &g  �<    0                   Kg  �<         jg  `B    R                   �g  `B         �g  ��                         �g  0B    0                   �g  0B         h  �i	         Bh  �l	         Xh  S                        zh  �l	         �h  �l	         �h   m	         �h  @p	         �h   S                        i  @p	         !i  p	         7i  `�                         Zi  �x                        }i  ��                         �i  �x                    .text   �                       .data                           .bss    P                            �i  @                               �i  h                        j  H                        5j  t                        [j  d                         �j  �                        �j  l                        �j  �                    .rdata  �     "                     �j  �i	    +                   &k  �                          Zk  �                         �k  �l	    H                    �k  �                          �k  �                         �k  �l	    0                     l  �                         l  �                         :l   m	                       ml  �                          �l  �                         �l  @p	    H                    �l  �                          m  �                         +m  p	    0                    Gm  �                         dm  �                         �m  ��                          �m   �         �m   �               *n   �         bn   �         �n   �         �n   �         o   �         Ho   �         �o   �         �o   �         �o   �         $p  0�         Hp  0�         |p  0�         �p  0�         �p  0�         q  0�         >q  0�         mq  0�         �q  0�         �q  0�         r  0�         %r  P�         Nr  P�         �r  P�         �r  P�         �r  P�         (s  P�         ]s  P�         �s  P�         �s  P�          t  P�         4t  P�         ]t  @�         �t  @�         �t  �>         �t  �<         u  �?         ;u  0G         mu  0D         �u  �H         �u  �L         v   J         >v  �M         tv  C	         �v  ��     X                   �v  C	         �v  px         �v  px         w  py         ;w  py         _w  pz         �w  pz         �w  �B	         �w   �     X                   �w  �B	         x        0x         1x  0x         Tx  0y         xx  0y         �x  0z         �x  0z         �x  �B	         y  @x         )y  @y         My  @z         vy  �B	         �y   x         �y   y         �y   z         �y  ��         Fz  p�         �z  �x         �z  �     X   
                �z  �x         	{  �x         +{  �y         N{  ��     X   
                u{  �y         �{  �y         �{  �z         �{  `�     X   
                |  �z         7|  �z         _|  0�         �|  `�         �|  �W          }  �W          2}  �E         q}   �         �}  �W          �}  `�         e~  �         �~   M         '  0?         e  �@         �  Ж         �  `=         �  Ц         c�  PD         ��  �F         ր  @�         '�  PG         e�  �H         ��  ��         �  PH         �  �I         P�   �         ��  �G         �   O               +�  @K         o�  ��         Ã   J         �  �M         G�  �         �  �?         ��   A         �   �          �  0�         I�  �M         ��  PL         ��  P         ��  Э         s�  `�         ��  �L         �  �>         %�   @         `�   >         ��  �         �  ��         �  �<         R�  0I         ��  ��         ��   �         �   �                         �  t                        #�   �     !                    O�  �|     8                   {�  p�                         ��   ~                        ��  ��     "                    މ  @|     8                   �  @�                         '�  �}                        C�  @�     "                    p�   |     8                   ��   �                         ��  �}                        Պ   �                         ��  �z                        #�        ��                         K�   {                        s�  ��     "                    ��   }                        ͋   �                         �  pz                        �  ��                         C�   {                        k�  @�     "                    ��   }                        Ō  @�                         �  �z                        �  ��                         8�  @{                        _�  ��     !                    ��  @}                        ��   �     X   
                Ӎ  ��     X   
                �  ��     X   
                �  P�     X   
                =�  0�     X   
                e�  ��     X   
                ��   �     X   
                ��  ��     X   
            .text   �                       .data                           .bss    P                            �  ��    �                    ,�  	                                r�  �                         ��   �                         �  	                          �  �                         S�  0�                         }�  	                          ��  �                         Ӑ  P�                         �   	                          2�                           b�  @�                         ��  $	                          ��                           �  �>                         �  (	                          W�                           ��  �<                         ƒ  ,	                          ��  (                         6�  �?                         l�  0	                          ��  4                         ړ  0G                         �  4	                          K�  @                         ��  0D                         ��  8	                          ��  L                               .�  �H                         e�  <	                          ��  X                         Օ  �L                         �  @	                          P�  d                         ��   J                         ˖  D	                          	�  p                         G�  �M                         ��  H	                          ��  |                         ��  C	                        �  L	                          :�  �                         Y�  px                        ��  P	                          ��  �                         ֘  py                         �  T	                          +�  �                         V�  pz                        ��  X	                          ��  �                         �  �B	                        �  \	                          "�  �                         A�  0x                              j�  `	                          ��  �                         ��  0y                        �  d	                          �  �                         >�  0z                        m�  h	                          ��  �                         ͛  �B	    $                    �  l	                          
�  �                         )�  @x    $                    R�  t	                          |�  �                         ��  @y    $                    М  |	                          ��                            &�  @z    $                    U�  �	                          ��                           ��  �B	    $                    ӝ  �	                          �                           �   x    $                    :�  �	                          d�  $                         ��   y    $                    ��  �	                                �  0                         �   z    $                    =�  �	                          m�  <                         ��  ��    -                     �  �	                          :�  H                         ��  p�    �                     �  �	                          H�  T                         ��  �x                        С  �	                          ��  `                         "�  �x    $                    J�  �	                          s�  l                         ��  �y                        Ţ  �	                          �  x                         �  �y    $                    B�  �	                          l�  �                         ��  �z                        ģ  �	                          �  �                         "�  �z    $                    P�  �	                          �  �                         ��  0�                              ��  �	                          ;�  �                         ��  `�    [                    إ  �	                          /�  �                         ��  �E    0                   ˦  �	                          �  �                         W�   �    3                    ��  �	                          �  �                         X�  `�    �                    �  �	                          q�  �                         ��  �    K                    ��  �	                          �  �                         ��   M    o                    ֫  
                          !�  �                         l�  0?                        ��  
                          ��  �                         :�  �@                        |�  
                          ��                           �  Ж    _                    ;�  
                                u�                           ��  `=    �                    �  $
                          8�                            }�  Ц    F                    ԯ  0
                          ,�  ,                         ��  PD    *                   Ȱ  8
                          �  8                         R�  �F    |                    ��  H
                          ɱ  D                         �  @�    �                    \�  X
                          ��  P                         �  PG    u                    P�  d
                          ��  \                         ڳ  �H    u                    �  l
                          _�  h                         ��  ��    n                    �  t
                          ;�  t                         ��  PH    5                    õ  �
                          ��  �                               ;�  �I    5                    u�  �
                          ��  �                         �   �    �                     K�  �
                          ��  �                         �  �G    �                    R�  �
                          ��  �                         ޸   O    	                   &�  �
                          o�  �                         ��  @K    	                   �  �
                          M�  �                         ��  ��    <                    �  �
                          M�  �                         ��   J                       �  �
                          ;�  �                         ��  �M                       ̼  �
                          �  �                         \�  �    �                    ��  �
                          ٽ  �                         �  �?    ,                          R�  �
                          ��  �                         Ⱦ   A    ,                    �  �
                          ;�                           u�   �    �                    ��  �
                          ��                           7�  0�    /                    f�                            ��                           ��  �M    ,                    �                            G�  (                         ��  PL    ,                    ��                            	�  4                         J�  P    ,                    ��  $                          ��  @                         	�  Э    2                   ��  ,                          �  L                         ��  `�    p                    ��  @                          �  X                         >�  �L    w                    ��  H                          ��        d                         �  �>    �                    ^�  P                          ��  p                         ��   @                        '�  X                          i�  |                         ��   >    q                    ��  `                           �  �                         [�  �    �                    ��  p                          �  �                         \�  ��    _                    ��  |                          ��  �                         �  �<    a                    I�  �                          ��  �                         ��  0I    �                    �  �                          X�  �                         ��  ��    k                    ��  �                          ��  �                         +�   �    �                    d�  �                          ��  �                         ��  �#                                ��  �#                          �  �W                          >�  �W                          e�  �W                          ��  ��                          ��  �          ��  �M                         �  �R                        !�  �           @�   M                        d�  `           ��   J                        ��  �           ��  0J                        �  �S                        S�              u�   N                        ��  �S                        �  @           8�  @N                        ��  0S                        ��              ��  �M                        J�  �          k�  �M                        ��  �          ��  �M                        ��  �R                        ��   !          �  M                        :�  �           ^�  @J                        ��  �           ��  PJ                               ��  �S                        )�  0           K�  0N                        ��  �S                        ��  P           �  PN                        `�  @S                        ��             ��  �M                         �  �          A�  �M                        f�  Љ         ��  �]     .text   �                       .data                           .bss    P                            ��  ��    �  �                 ��  �     Z                    �  �                         J�  Љ    �  M                 ~�       |                    ��  �                         ��  �]    Y                   �  �     ,                    �  �                         ;�  �                           b�                             ��  P                           ��  0                           ��  �                           �  �                 !                -�  �                          T�   !                          y�  �                           ��                              ��  @                           ��                              �  `                           A�  �                           k�  �                          ��  �                           ��                             �  �!         ��  �#         2�  �"         ��             ]�   !         ��  �"         8�   -         ��  �6         @�            ��  �         ��  �         �  `&         ��  @(         J�  `'         ��  �$         u�  �%         	�  @'         P�  �2         ��  �9         X�             ��  �         ��  �8         o�  �5         ��  �         6�  `         ��  �         ��  �         $�  ��         `�  0�         ��  p�         ��  �          �  p�         F�  ��         �  �        "        ��  ��         ��  ��         )�  0�          a�  ��         ��  P�         ��  p�          �  P�         D�  0�         ~�  ��          ��  0�         ��  �         +�  P�          d�  �         ��  ��         ��  ��          �  ��         K�  ��         ��  �          ��  ��         ��  P�         1�  �          i�  P�         ��  p�         ��  ��          �  p�         L�  ��         ��  �          ��  ��         �  0�         G�  �          ��  0�         ��  ��         �  е          A�  ��         ��  p�         ��  ��          ��  p�         <�  �         u�  ��         ��  P�         ��  p�          �  P�         U�  P�         ��  p�         ��  0�         �  �         ;�  �          r�  �         ��  ��         ��  ��         �  ��         V�  ��         ��  ��         ��  ��         �  ��         F�  P�         ��  ��#               ��  p�         ��  ��         4�   1         ��  @+         ]�  �r                        ��  �r         ��  ��    �                  8�  ��         ��  0�    (                  0�  0�         ��  ��                        �  ��         ��  ��                        ��  ��         Y�  0�    �                   ��  0�         O�  p�    �                   ��  p�         E�  @�    J                  ��  @�         W�  �    J                  ��  �         i�  �    �                  ��  �         {�  p�    �                    p�         �  P�    �                   �  P�         Y `�    �                   � `�         % ��                      � ��           �                      �  �          p�                        c p�         � ��                        ! ��         } ��    $                          � ��         o ��                        � ��         a ��    �                   ��         � п    �                  n	 п         
 ��    �                  �
 ��         � p�    �                  \ p�          0�    G                  � 0�         w ��    G                  ) ��         � `           �l                        $ �f          \ ��          � �d          � ��           @k          @  �          ~ �j          � ��          � �h          3 ��          l �i          � ��          � �e           ��          N @g          �  �          � @e          �  �          , @l          j  �          � �k          � ��          $ @i          ]  �          � @j          �  �           @f          @  �          x ��                         � %      �g          � ��           @h          D  �      .text   �                       .data                           .bss    P                            |      ,                    � �                          %  	                         z �!    n                     �                          � 	                         J �#    n                    � �                          � 	                         ) �"    n                    � �                          d $	                                n                    � �                          7 0	                         �  !    n                    l  �                          ! <	                         �! �"                        �! �                          =" H	                         �"  -    �                    # �                          �# T	     &                          I$ �6    n                    �$ �                          J% `	                         �%                          & �                          Z& l	                         �& �    #                    �& �                          K' x	                         �' �    ,                    �'                            I( �	                         �( `&    n                    8)                           �) �	                         n* @(    n                    +                           �+ �	                         M, `'    n                    �,                           �- �	                         &. �$    n                    �.                            [/ �	                         �/ �%    n                    �0 (                          +1 �	                         �1 @'        '                      2 0                          a2 �	                         �2 �2    �                    C3 4                          �3 �	                         m4 �9    n                    �4 @                          n5 �	                         �5                           66 H                          ~6 �	                         �6 �    #                    7 L                          o7 �	                         �7 �8                        R8 T     *                    �8 
                         p9 �5                       �9 �     *                    w: 
                     .rdata  �     �   ,                 �: �    �                    K; �     !                    �;  
                         �; `    �                    =< �     !                    �< ,
                         �< �    �            (              D= �     $                    �= 8
                         > �    �                    [>      $                    �> D
                         �> ��    4                    5? <                          x? P
                         �? 0�    4                    �? D                          @@ \
                         �@ p�    0                    �@ L                          A h
                         BA ��    >                    �A T                          �A t
                         B ��    >                    @B \                          �B �
                         �B P�    0                    �B d                          ?C �
                         C 0�    >                    �C l                           D �
                         AD �    >                    �D t                          )      �D �
                         E ��    >                    CE |                          �E �
                         �E ��    >                    F �                          FF �
                         �F P�    <                    �F �                          G �
                         FG p�    <                    �G �                          �G �
                         H ��    `                    JH �                          �H �
                         �H 0�    `                    I �                          aI �
                         �I ��    `                    �I �                          2J �
                         xJ p�    `                    �J �                          K                          IK �    F                    �K �                          �K                          L �� *         F                    GL �                          �L                          �L P�    G                    M �                         DM (                         �M P�    F                    �M �                          N 4                         EN p�    F                    �N �                          �N @                         O 0�    F                    GO �                          �O L                         �O �    G                    P �                         FP X                         �P ��    8                    �P                           Q d                         DQ ��    F                    �Q                           �Q p                         R ��    8                    ER                           �R |                         �R ��    D                    S       +                          DS �                         �S ��    D                    �S $                          T �                         CT ��    h                    �T ,                          �T �                         U ��    h                    YU 4                          �U �                         �U P�    h                    *V <                          pV �                         �V ��    h                    �V D                          AW �                         �W p�    O                    �W L                         X �                         CX ��    O                    �X \                         �X �                         �X  1    �                   �Y l     9                    @Z �                         �Z @+    �                   v[ �     9                    \ �             ,                  �\ �                         �\                          ] �     <                   �]                         ^ $     L                   �^                         _ p                         v_ $                        �_ t                         V` 0                        �` x     !                   Ea <                        �a �     !                   Cb H                        �b �     H                   Oc T                        �c      H                   id `                        �d P     ^                   �e l                        f �     ^                   �f x                        *g      !                   �g �                        �g 4     !                   hh �                        �h X     +                   Mi �                    -          �i �     +                   Cj �                        �j �                         !k �                        �k �                         �k �                        Jl �                         �l �                        Dm �                         �m �                        >n �                         �n �                        �o �                         Tp �                        q �     4                   �q �                        �r      5                   Rs                         t <     /                   �t                         |u l     /                   /v                          �v `    ;	  q                 w �     �                    Ew ,                         ww �f     8                    �w ��     5                     �w �d     8                    3x .      ��     4                     qx @k     8                    �x  �     ;                     �x �j     8                    @y ��     ;                     �y �h     8                    �y ��     6                     z �i     8                    Ez ��     6                     �z �e     8                    �z ��     5                     { @g     8                    B{  �     5                     �{ @e     8                    �{  �     4                     �{ @l     8                    B|  �     ;                     �| �k     8                    �| ��     ;                     } @i     8                    Q}  �     6                     �} @j     8                    �}  �     6                     ~ @f     8                    P~  �     5                     �~ �g     8                    �~ ��     5                      @h     8                    L  �     /      5                     � �     H                    � �     8                    � �     h                    M� �     h                    �� ��     0                    Ҁ P�     0                    � �     8                    Q� ��     H                    �� p�     8                    ΁ ��     h                    � е     h                    X� �     0                    �� ��     0                    ؂ p�     8                    � 0�     P   	                 V� �     P   	                 �� ��                        �� ��                          �� @s                        ԃ @s         � p�                        �� p�         � ��                        $� ��         7�  �                        N�  �         _� P�    +                   z� P�         �� ��    +                   �� ��         ф ��         0                     � ��         �� ��                        � ��         3�  s                       N�  s         c� ps                       ~� ps         �� `x    $                   �� `x         Å �d                       	� �d         I� �d                       �� �d         ц  e                       �  e         � �d                       3� �d         Q� Pb                        l� Pb         �� �d                       �� �d         �� �                          ۇ Ѐ                       � Ѐ         �� ��                       � ��         � @�                        $� @�         3� ��                        F� ��         S� ��                        i� ��         y�  �    
                    ��  �         �� ��                        �� ��         �� 0�                 1             Ո 0�         � @�                        �� @�         � `�    
                     � `�         /� 0�                        C� 0�         Q� ��                        g� ��         w� ��                        �� ��         �� ��                        �� ��         ˉ p�                        �� p�         � ��                         � ��         � ��    %                   � ��         )� ��                        >� ��         M�  �                        a�  �         o� @�    l                   �� @�         �� �h    .                    �� �h         �� ��                       ͊ ��         ي �m                       �� �m         � P�                        � P�         %� ��                        9� ��         G� ��                        e� ��         }� ��    �   2                      �� ��         �� ��                       �� ��         ы ��    0                   � ��         �� ��    B                   � ��         � ��    l                   6� ��         I� 0�                       b� 0�         u� ��    0                   �� ��         �� @�    0                    �� @�         Ō  �    r                   �  �         � ��                       %� ��         A� ��    0                   b� ��         }� ��                       �� ��         �� �    s                   ֍ �         � ��                       � ��         -� ��    0                   M� ��         g� ��    0                    �� ��         �� ��    r                   Î ��         � `�                       	� `�         )� ��    0                   N� ��         m� p� 3         D                    �� p�         �� �    Z                   ҏ �         � p�                       � p�         5� ��    0                   Y� ��         w� ��    0                    �� ��         �� ��    Q                   ϐ ��         �  �    �                   ��  �         � ��    �                   3� ��         K� �    b                   d� �         w� ��    �                   �� ��         �� ��    ~                   Ñ ��         ّ �b                        �� �b         � pb                        E� pb         e�  g                       ��  g         ��  �                        Ò  �         ߒ �    	                    � �         � 0g                        ?� 0g         [� @g                        � @g         �� Pg                        ̓ Pg       4        �� g                        � g         -�  h    {                   R�  h         q� �x    ^                  �� �x         �� �b    /                   �� �b         є Ps                       � Ps         �� �h    .                   
� �h         � 0j                        +� 0j         9� ��    (                   I� ��         S� i                        g� i         u� pr    2                   �� pr         �� �f    $                   �� �f         �� �h    0                   ʕ �h         ו `f    >                   � `f         � 0i                       � 0i         � �i    L                   *� �i         9� Pi    4                   q� Pi         �� �i    E                   ޖ �i         � `e    |                   4� `e         O� po    &                   e� po5               u� p�    ,                   �� p�         ��  r    C                   ��  r         �� �o    =                   � �o         %� Pw    K                   >� Pw         Q� �t                       �� �t         ɘ �o    !                   � �o         9� �e    b                   ]� �e         {� �m    �                   �� �m         �� P�                        ˙ P�         � o    C                   � o         � �m    (                   0� �m         A� �    (                   S� �         _� `o                       �� `o         �� Pp    m                  Ț Pp         ۚ �o                       +� �o         u� �q    L                   �� �q         ��  p    0                   ��  p         ϛ �q                       � �q         ��  x    >               6          �  x         #� �b    W                   G� �b         e� �                       u� �         � �|                       �� �|         �� 0~                       �� 0~         ��  {                       ՜  {         �  �                        ��  �         � �|                        '� �|         9� �}    %                   K� �}         W� Pz    %                   i� Pz         u� Pf                       �� Pf         Ý �f                       � �f         � �f                       ,� �f         K�  g    
                    j�  g         �� �g    l                   �� �g         Þ �w    q                   ٞ �w         �  e    ?                   �  e         � pk    �                   5� pk         G�  �                       Z�  �         g�  l    �      7                   ��  l         �� �j    �                   �� �j         �� �                       � �         � Pj    (                   � Pj         -� Ё    (                   ?� Ё         K� �l                       v� �l         �� �l         �� �l                       ɠ �l         ٠ �r    _                   � �r         �� �r                       � �r         #� �y    W                   ;� �y         M�  �    Z                   ]�  �         g� `g    (                   �� `g         ��  {    F                   ��  {         ɡ P~    F                   ܡ P~         � �n    _                   � �n         � @�                       &� @�         3� P�	    �                   p� P�	         �� P�	    z                   � P�	         � ��	    l                   R� ��	    8           ��  c    k                   �  c         S�  �    "                   ��  �         Ѥ �|    "                   � �|         O� d    x                   �� d         ե �~    F                   � �~         � p{    F                    � p{         5� �~    W                   J� �~         Y� �{    W                   n� �{         }� ��    9                   �� ��         �� P    W                   �� P         צ  |    W                   �  |         	� ��    "                   (� ��         A� P}    "                   `� P}         y� �c    x                   �� �c         ��  ~    &                   �  ~         -� �z    &                   G� �z         [� 0u    �                  v� 0u         �� �v                       �� �v         �� �v    R                   ب9       �v         � �t    ;                   	� �t         �  t                       ^�  t         �� 0t    #                   ک 0t         � �s    A                   U� �s         �� `t                       Ҫ `t         �  t                       R�  t         �� �t    #                   � �t         1� �t                       t� �t         �� �s                       �� �s         C� �}    C                   \� �}         o� �z    C                   �� �z         �� �    &                   ȭ �         � �|    &                   � �|         C� P�    "                   c� P�         }�  }    "                   ��  }         �� ��    
                    �� ��         3� ��    
                    u� ��         �� ��         ӯ  �         �� `V                         � PV   :                            =� pV                     .text   �                       .data                           .bss    P                            P� P                         h� 8                        �� T                         �� D                        �� X                         ǰ P                        ް \                         �� \                        � `                         *� h                    .rdata  �                         B� d                         ^� t                        z� l                         �� �                        ı t                         ޱ �                        �� x                         � �                        6� |                         R� �                        n� �                         �� �                        �� �        ;                       ² �                        ޲ �                         %� �                        l� �                         �� �                        �� �                         � �                        B� �                         g� �                        �� �                         �� �                        Ĵ �                         �                         �� �                         �                          � �                         1�                         B� �                         X� (                        n� �                         �� 4                        �� �                         �� @                        ĵ �                         ٵ L                        � �                         � X                        � �                <               1� d                        F� �                         ^� p                        v� �                         �� |                        �� �                         �� �                        ̶ �                         � �                        �� �                         � �                        ,� �                         E� �                        ^� �                         t� �                        �� �                         �� �                        �� �                         �� �                        Է �                         � �                         � �                         � �                        *� �                         B� �                        Z� �                         p�                          �� �                       =        ��                         ��                          ĸ                         ܸ                          � $                        �                          � 0                        2�                          Q� <                        p�                          �� H                        �� ,                         �� T                        Թ 0                         � `                        � <                         � l                        0� H                         J� x                        d� X                         ~� �                        �� \                         �� �                        ʺ h                         � �                        �� l                         � �                        >� |                         a� �>                              �� �                         �� �                        Ȼ �                         � �                        � �                         *� �                        L� �                         n� �                        �� �                         �� �                        Ҽ �                         � �                        � �                         7�                         ^� �                         ��                         �� �                         ҽ                          �� �                         � ,                        @� �                         f� 8                        �� �                         �� D                        ؾ �                         �� P                        "� �                         E� \     ?                         h� �                         �� h                        ��                          �� t                        ؿ                          �� �                        �                           0� �                        J� 0                         f� �                        �� @                         �� �                        �� L                         �� �                        
� P                         1� �                        X� T                         z� �                        �� X                         �� �                        �� \                         � �                        (� `                         K� �                        n� d                         �� �                        �� h                         ��            @                   � l                         8�                         X� p                         ~�                         �� x                         �� (                        �� �                         �� 4                        � �                         +� @                        B� �                         V� L                        j� �                         � X                        �� �                         �� d                        �� �                         �� p                        �� �                         �� |                        � �                         � �                        2� �                         F� �                        Z� �                         l� �                        ~� �                         �� �                  A            �� �                         �� �                        �� �                         � �                        F�                          �� �                        ��                          �� �                        � $                         � �                        0� ,                         A� �                        R� 4                         j�                          �� <                         ��                         �� H                         �                         ,� P                         l� $                        �� T                         �� 0                        $� \                         I� <                        n� l                         �� H                        �� x                         �� T                        ��B       �                         	� `                        $� �                         <� l                        T� �                         g� x                        z� �                         �� �                        �� �                         �� �                        � �                         W� �                        �� �                         �� �                        �� �                         �� �                        � �                         ,� �                        F� �                         ^� �                        v� �                         �� �                        �� �                         �� �                        �� �                         �� �                        � �                         � �                        2� �   C                            I�                         `�                          y�                         ��                          ��                          ��                          �� ,                        ��                          �� 8                        � $                         ;� D                        f� (                         �� P                        �� ,                         �� \                        �� 0                         � h                        >� 4                         b� t                        �� @                         �� �                        �� H                        �� �                        �� d                         	� �                        "� t                         6� �                        J� x        D                       e� �                        �� �                         �� �                        �� �                         �� �                         � �                         � �                        0� �                         C� �                        V� �                         �� �                        �� �l    �                    �� �                          �� �                         
� �                         !�                         8� �                         O�                         f� �                         |�                         �� �                         �� (                        �� �                         �� 4                        �� �                         � @                        0� �                         D� L               E               X�                          l� X                        ��                          �� d                        ��                          �� p                        ��      %                   � |                        V� D     $                   �� �                        �� h                        
� �                        F� �                         �� �                        � �                         ]� �                        �� �                         �� �                        &� �                         m� �                        �� �                         �� �                        �� �                         � �                        $� �                         :� �                        P� �                         f� �                      F        |� �                         ��                          �� �                         ��                         �� �                         �                          � �                         @� $                        `� �                         �� 0                        �� �                         �� <                        .�                           I� H                        d�                          � T                        ��      ,                   �� `                        �� <                         �� l                        
� D                         (� x                        F� L                         a� �                        |� \                         �� �                         � `                         B� �                        �� hG                               �� �                        � x                         J� �                        �� |                         �� �                        � �                         k� �                        �� �                         � �                        H� �                         �� �                        �� �                         �� �                        � �                         0� �                        J� �                         x�                         �� �                         ��                         � �                         #�                          D� �                         e� ,                        �� �                         �� 8                        
� �                         M� D                        �� ��    H      �                    �� �                          �� P                         
�  �    �                    :� �                          k� \                         ��  �                        ��  �                          �� ��                        )� ��         T� p�                        �� p�         �� p�                        �� p�         � �                        ?� �         j�  �    +                   ��  �         �� ��    +                   � ��         D� 0�                        w� 0�         �� ��                        �� ��         � ��    '                   C� ��         r�  �    '                   ��  �         �� ��    %                    � ��         :� p�    '                   �� p�         �� @�    '                   Z� @�         �� ��    '                   �� I      ��         ,� ��    '                   j� ��         �� ��                        �� ��         � 0�                       <� 0�         l� �                          �� ��                       �� ��         �� `�                       &� `�         J� �                        y� �         �� ��                        �� ��         �� ��                        &� ��         P� ��    
                    ~� ��         �� ��                        �� ��          �  �                        .�  �         V� ��                        �� ��         �� 0�    
                    �� 0�         
�  �                        8�  �         `� ��                        �� ��         �� `�                        �� `�         � P�                        J� P�         v� @�                        �� @�    J           �� ��                        �� ��         � ��    &                   J� ��         p� P�                        �� P�         �� ��                        �� ��         � �    o                   O� �         z� �    .                    �� �         �� ��                       � ��         (� ��                       Z� ��         ��  �                        ��  �         �� ��                        � ��         4� ��                        l� ��         �� ��    �                    �� ��         �� ��                       /� ��         \� ��    0                   �� ��         �� ��    J                    �� ��         � ��    �                    C� ��         p�  �                       ��  �         �� `�    0                   � `�         0� 0�    1                    `�K       0�         ��  �    G                    ��  �         �� p�                       9� p�         p� ��    0                   �� ��         �� ��                       � ��         L� @�    S                    �� @�         �� ��                       �� ��         .� �    0                   h� �         �� ��    1                    �� ��         � ��    Y                    F� ��         �� 0�                       �� 0�         �� ��    0                   ;� ��         t� @�    D                    �� @�         ��  �    N                    '�  �         `� P�                       �� P�         �� ��    0                   � ��         P� `�    1                    �� `�         �� ��    h                    �� ��         &�  �    �                   ]�  �         �� ��               L             �� ��         ��  �    �                   -   �         Z  P�    �                   �  P�         �  P�    �                   �  P�         $ ��                        b ��         � ��                        � ��          �                       K �         � ��                        � ��         � ��    	                    . ��         d  �                        �  �         � 0�                         0�         L @�                        � @�         �  �                          �         D �    �                   � �         � ��    K                  � ��           �    /                   P  �         �  �                       �  �         � ��    .                    ��         . `�                        \ `�         � @�        M                      � @�         � P�    )                    P�         ( �    6                   W �         � ��    1                   � ��         � ��    (                    	 ��         &	 P�    ?                   Q	 P�         v	 `�                       �	 `�         �	 �    L                   �	 �         $
 ��    7                   w
 ��         �
 ��    I                    ��         j @�    �                   � @�         � ��    &                   
 ��         4  �    ,                   ^  �         � ��    C                   � ��         � 0�    @                   3 0�         � p�    K                   � p�         � ��                       < ��         � p�    $                   � p�         6 ��    c                   t ��         � 0� N         �                   � 0�         
  �                        J  �         � ��    D                   � ��         �  �    (                     �         D ��    (                   p ��         � ��                       � ��          ��    �                  M ��         z �                       � �         J p�    L                   � p�         � ��    0                   � ��          `�                       B `�         p @�    >                   � @�         � 0�    f                    0�         > ��                        n ��         � 0�                        � 0�         � @�                       4 @�         p p�    7                   � p�         � ��    7                   � ��          ��    5                   : ��       O        b  �    5                   �  �         � ��    =                   � ��          `�    =                   9 `�         ` ��                       � ��         � ��                        ��         H ��    
                    � ��         � ��                       � ��         $ ��    q                   T ��         ~  �    ?                   �  �         � ��    �                    ��         F ��                       t ��         � 0�    �                   � 0�           ��    �                   2 ��         ^ ��                       � ��         � ��    (                   	 ��         4 ��    (                   ` ��         � ��                       � ��         
  �         <  �                       l  �         � `�    _        P                 � `�         � P�                        P�         H  �    S                   z  �         � ��    V                   � ��         � `�    (                   0  `�         f  `�    F                   �  `�         �  ��    F                   �  ��         !  �    _                   E!  �         r! ��                       �! ��         �! p�	    �                   " p�	         <" ��	    �                   w" ��	         �" �	    l                   �" �	         # ��    m                   �# ��         $ ��    "                   u$ ��         �$ P�    "                   %% P�         z% ��    �                   �% ��         0& 0�    G                   d& 0�         �& ��    G                   �& ��         �& ��    Y                   $' ��         N'  �    Q      Y                   ~'  �         �' ��    9                   �' ��         ( ��    Y                   9( ��         h( `�    Y                   �( `�         �( 0�    "                   ) 0�         4) ��    "                   k) ��         �) �    �                   �) �         R* p�    &                   �* p�         �* ��    &                   �* ��         + @�    �                  C+ @�         r+ ��                       �+ ��         �+ �    R                   , �         B,  �    ;                   v,  �         �,  �                        -  �         V-  �    &                   �-  �         
. ��    G                   e. ��         �. P�    !                   / P�         p/ ��    !                   �/ ��         &0 ��    ,                   �0 ��         �0 R      ��    !                   \1 ��         �1 P�    !                   2 P�         ~2  �    C                   �2  �         �2 ��    C                   3 ��         63 @�    $                   {3 @�         �3 ��    $                   �3 ��         >4  �    "                   v4  �         �4 ��    "                   �4 ��         5 ��    
                    m5 ��         �5 ��    
                    6 ��         t6 0V                         �6  V                         �6 @V                     .text   �                       .data                           .bss    P                            7 �                         G7 h                        y7 �                         �7 t                        �7 �                         8 �                        ?8 �                         s8 �     S                         �8 �                         �8 �                    .rdata  �     �                    9 �                         A9 �                        w9                          �9 �                        �9                          ): �                        ]:                          �: �                        �:                          ; �                        ;;                          q; �                        �;                          �; �                        <                           v< �                        �< $                         <=                         �= (                         �=                         > ,                         \>                         �> 0                         �> (                        ? 4          T                     >? 4                        u? 8                         �? @                        �? <                         �? L                        !@ @                         Q@ X                        �@ D                         �@ d                        �@ H                         A p                        ?A L                         nA |                        �A P                         �A �                        �A T                         .B �                        ]B X                         �B �                        �B \                         �B �                        !C `                         PC �                        C d                         �C �                        �C h                         D �                        GD l                  U             zD �                        �D p                         �D �                        E t                         9E �                        eE x                         �E                          �E �                         �E                         F �                         NF                         }F �                         �F $                        �F �                         G 0                        CG �                         qG <                        �G �                         �G H                        H �                         5H T                        eH �                         �H `                        �H �                         �H l                        5I �                         hI x                        �I �                         V      �I �                        J �                         5J �                        gJ �                         �J �                        �J �                         �J �                        /K �                         dK �                        �K �                         �K �                        �K �                         0L �                        aL �                         �L �                        �L �                         M �                        WM �                         �M �                        �M                           	N �                        CN                          N                         �N                          �N                         5O                          pO                          �O                          �O ,  W                            P                          ^P 8                        �P $                         �P D                        #Q (                         cQ P                        �Q 4                         �Q \                        R 8                         _R h                        �R <                         �R t                        !S @                         `S �                        �S L                         �S �                        T P                         OT �                        �T T                         �T �                        �T \                         /U �                        iU h                         �U �                        �U t                         V �                        =V �                         tV �      X                        �V �                         �V �                        )W �                         hW �                        �W �                         �W �                        X �                         \X                         �X �                         �X                         Y �                         PY                         �Y �                         �Y (                        Z �                         UZ 4                        �Z �                         �Z @                        [ �                         Q[ L                        �[ �                         �[ X                        �[ �                         0\ d                        g\ �                         �\ p                        �\ �                         �\ |             Y                 %] �                         T] �                        �] �                         �] �                        �] �                         ^ �                        7^                          g^ �                        �^                          �^ �                        �^                           _ �                        M_ $                         y_ �                        �_ 0                         �_ �                        ` 4                         3` �                        c` <                         �` �                        a H                         ba                          �a T                         �a                         1b d                         bb                         �b l                         �b $                    Z          �b t                         c 0                        Mc |                         �c <                        �c �                         -d H                        ad �                         �d T                        e �                         ne `                        �e �                         f l                        Cf �                         vf x                        �f �                         �f �                        +g �                         ag �                        �g �                         �g �                        �g �                         (h �                        Uh �                         �h �                        �h �                         i �                        Ii �                         �i �                        !j [      �                         Xj �                        �j                           �j �                        �j                          *k �                        _k                          �k �                        �k                           l                         =l $                         nl                         �l ,                         �l                          m 4                         Dm ,                        �m 8                         �m 8                        �m @                         n D                        3n H                         bn P                        �n P                         �n \                        �n X                         o h                        Ko `                         yo t                        �o h     \                          �o �                        #p l                         ap �                        �p p                         �p �                        q t                         Oq �                        �q �                         �q �                        �q �                        %r �                        ]r �                         �r �                        �r �                         �r �                        #s �                         Ys �                        �s �                         �s �                        �s �                         6t �                        wt �                         �t                         �t �                         u                         5u �                         {u                         �u  �    �    ]                      �u �                          2v (                         kv                          �v 4                        �v                          �v @                        /w                          _w L                        �w                          �w X                        �w (                          x d                        Kx 4                         �x p                        �x 8                         �x |                        #y @                         Ry �                        �y H                         �y �                        �y T                         z �                        Gz X     &                   �z �                        �z �     %                   �z �                        ;{ �                        w{ �                 ^             �{ �                         6| �                        �| �                         } �                        q} �                         �} �                        )~ �                         �~ �                        �~ �                                                   Q �                         �                         �                           �                         �                           N� $                        �                           �� 0                        �                           � <                        O� $                          �� H                        �� ,                          � T                        +� 4                          c� `                        �� <                          �� l                        _      Y� L                          �� x                        �� T                          � �                        %� \      ,                   [� �                        �� �                          Ȅ �                        �� �                          8� �                        q� �                          �� �                        ۅ �                          8� �                        �� �                          � �                        Q� �                          �� �                        	� �                          h� �                        ǈ �                          &� �                        �� �                          �� �                        e� �                          Ċ                         #� �                          ��                         �� �   `                             '�                          Y� �                          �� ,                        �� �                          � 8                        I� �                          �� D                        Ս !                         � P                        G� !                         �� \                        �� !                         � h                        q� !                         Ώ t                        +�  U                        L�  U                          g� 0U                        �� 0U         �� ��         �� ��     `                   ѐ ��         � ��         ��  �     �                   � @R                        >� ��         Q� �         l� �         �� ��         �� p�         �� ��         ȑ U                       � U       a        � �T                       >� �T         `� PS         �� �R         �� �         �� �         ɒ ��         ޒ ��         � и         � p�     �                   0� и         N�  �                         h� pr                        ��  �                         �� `}     8                   ��  �                         ؓ �{     8                    � �                         � �}                        .� @�                         M� @t                    .text   �                       .data                           .bss    P                            l� !                         �� �                        ��  !                         Ԕ �                        �� ��    <                    � $!                         +� �                         E� ��    6                    ^� 4!             b                  x� �                         �� �    6                    �� D!                         Օ �                         �� ��                        � T!                          *� �                         D� p�    >                    ]� \!                         w� �                         �� ��    >                    �� l!                         Ԗ �                         �� |!                         !� �                        L� �!                         u� �                        �� PS    �                    Ɨ �!                          � �                         � �R    �                    ?� �!                          g�                           �� �    [                    �� �!                                                    ܘ ��    C                    �� �!                      c          �                       .rdata  �                          /� и    �                    S� �!     &                    x� (                          ��  X                          �� 0"                          ٙ  "                          � �V                          � �V                          2� �V                          R� 0W                          s�  W                          �� �V                          �� �V                          Ӛ �V                          �  W                          � �V                          3� �V                          S� W                          s� �R                          ��  R         �� �         ϛ ��          � @�         � pR                        ;� @�         T� �         k� �         �� @R         �� �Q     .text   �                       .data                 d                .bss    P                            Ɯ �R                         � �!                          � 4                          4�  R                         X� �!                          }� @                          �� �                        ȝ  "                          � L                          � @�                        5� "                          U� X                          u� �    ~                    �� "                          �� d                          Ξ @R    ]                    �� "                          � p                          H� �Q    ]                    p� $"                          �� |                           ��                          L�                               ��              �� ��         � �     `                   7� ��         R� ��         �              >�         e           m� з         �� з         �� �V         Р @V         � �U         � �U         .� �U         P� pX         i� �W         �� @U         �� PV         ѡ Y         � �X         �  Z         +�  Y         O�  �         u�  �                         ��  t                    .text   �                       .data                           .bss    P                            �� ��                        Ԣ 4"                          �� �                          � ��    $                    9� 8"                          [� �                      .rdata  �     Q                     }� з    �                    �� @"     &                    ƣ �                          � �V    <                   � h"                          F� �                          t� @V                        �� l"                          ��f       �                          � �U    A                    
� p"                          3� �                          \� �U                        �� |"                          �� �                          ʥ �U    A                    � �"                          � �                          D� pX    [                    c� �"                          �� �                          �� �W    �                    Ȧ �"                          � �                          � @U    M                     >� �"                          i�  !                         �� PV    M                     �� �"                          � !                         � Y                         8� �"                          Z� !                         |� �X    1                     �� �"                          ͨ $!                         ��  Z  g        ;                    � �"                          =� 0!                         a�  Y    �                    �� �"                          �� <!                         �  �    �                    � �"                          :� H!                         L�                               ��              g� �v    	                    �� �v         ٪ �w    	                    � �w         K� �v                        �� �v         �� pu                        � pu         %� `u                        ^� `u         �� 0{    	                    ͬ 0{         � �{    	                    ?� �{         u�  {                        ��  {         � �y                        � �y         O� �y                        �� �y         �� �%	                       � �%	         �  �     h                   K� �)	       h                      }� �)	         �� ��     h                   ۯ `�    	                    � `�         ?� p�    	                    t� p�         �� p	                       ϰ p	         �� ��     H                   !� `�                        � `�         ױ ��                        :� ��         �� Щ                        ò Щ         �  �    "                    �  �         A� �@	                       �� �@	         ݳ @�     0                   .� �A	                       � �A	         ʴ ��     0                   � �?	                       k� �?	         �� ��     X   
                � !	                       ]� !	         >�              �� �%	    $                   � �%	         � P)	    $                   ?� P)	         k� �@	    $                   �� �@	         � �A	    $          i               X� �A	         �� @	    $                   ϸ @	         �� �?	    $                   E� �?	         �� � 	    $                   � � 	         9� 6	    (                   ]� 6	         {� `�     8                   �� �5	    0                   ú �5	         � �2	    (                   � �2	         !� �     8                   D� `2	    0                   g� `2	         �� P	    (                   �� P	         ֻ  	    0                   �  	         (� 0	    (                   S� 0	         x�  	    0                   ��  	         ȼ ��    &  	                � ��         4� 0B         v� �x    H                   �� �x         ޽ �z    H                   � �z         L� �{    H                   �� �{         �� @{    H                   �� @{         0� �v    H                 j        j� �v         �� Pw    H                   ڿ Pw         � �t    H                   G� �t         x�  w    H                   ��  w         �� �    H                   � �         D� `�    H                   t� `�         �� ��    H                   �� ��         �� �                       /� �         ^� ��	    �   
                �� ��	         �� 0T    o                   �� 0T         �� `�    L                   � `�         <�  �     h                   g� p�    L                   �� p�         �� ��    H                    � ��         C� Ь    H                   �� Ь         �� �    G                   �� �         )�  �    G                   Y�  �         �� 0u    #                   �� 0u         �� `v    #                   (� `v         [� �w    o                   �� �wk               �� @t    o                   �� @t         #� �u    o                   \� �u         �� �u    o                   �� �u         ��  u    #                   2�  u         c� t    #                   �� t         �� �s    #                   �� �s         /�  �    L                   Z�  �         � p�     h                   �� 0�    L                   �� 0�         �� ��    H                   C� ��         �� ��    H                   �� ��         � б    G                   B� б         l� �    G                   �� �         �� py    #                   �� py         2� �z    #                   k� �z         �� �{    o                   �� �{         �� �x    o                   5� �x         f� 0z    o                   �� 0z         �� �y    o                   � �y     l          >� @y    #                   u� @y         �� Px    #                   �� Px         �  x    #                   B�  x         r� �#	    �                   �� �#	         ��  "	    �                   �  "	         :� �$	    �                   �� �$	         �� �"	    �                   T� �"	         �� �%	                       �� �%	         � �'	    �                   A� �'	         p� �%	    �                   �� �%	         �� p(	    �                   4� p(	         �� �&	    �                   �� �&	         H� �)	                       z� �)	         �� �@	                       �� �@	         B� `@	                       �� `@	         �� �E    k                    W� �E         �� PE    k                    _� PE         �� �@	                       ?� �@	         �� �A	                       �� m      �A	         &� �A	                       w� �A	         �� Pm    ^                    '� Pm         �� �l    S                    	� �l         ��  B	                       ��  B	         "� �x    �  ,                �� �x         >� �"                         i� 0p    J  -                �� 0p         �� �"                         �� n                      � n         z� �m    ^                    � �m         ��  ;	    I                   ��  ;	         �� �     H                   �� :	    I                   
� :	         (� `:	    E                   d� `:	         �� p9	    E                   �� p9	         � �:	    G                   2� �:	         R� �9	    G                   x� �9	         ��  �    #                   ��  �         �� 0�    #                   (� 0�         T� ��    o             n            �� ��         �� �    o                   �� �         �� `�    o                   %� `�         L� �	    �                   {� �	         �� �	    �                   �� �	         �� `	    �                   V� `	         �� �	    �                   � �	         X� �	                       �� �	         �� �5                       !� �5         �� pQ                        ��  5                       _�  5         �� `?	                        � `?	         j� @?	                       �� @?	         � ��    #                   _� ��         �� ��    _                    2� ��         �� ��    _                    (� ��         ��  �    _                    "�  �         �� p�    _                    "� p�         �� @�    _                    � @�         �� �?	                       ��o       �?	         0� е    9                  �� е         6� @�    �                  �� @�         4� P�                      �� P�         R� �                      �� �         V� 0�                      �� 0�         ^� � 	                       �� � 	         � `�     X   
                f� ` 	                       �� ` 	         � � 	                       �� � 	         �� � 	                       u� � 	         ��  !	                       >�  !	         �� �5	    B                   �� �5	         �� �4	    B                   �� �4	         � @5	    B                   =� @5	         `� �4	    B                   �� �4	         �� �    #                   � �         f� @�    #                   �� @�         &� �    ,                    }� �         �� p�                       �� p�  p             � @6	    (                   >� @6	         \� ��                        �� ��         � ��                        X� ��         �� `	    �   
                �� `	         �� @�     8                   � �	    �   
                ?� �	         h� 	                       �� 	           P	                       p  P	         �  �	    (                   �  �	          p�         g p�         � 0    �                    0         h  Q                        � P    �                   � P         C 2	    B                   f 2	         � �1	    B                   � �1	         � �1	    6                   � �1	          @1	    6                   , @1	         K �                        � �         � P�                        � P�          �    #                   q      7 �         ] �2	    (                   � �2	         � @	    �                   � @	         � ��     8                    �	    �                   L �	         t  	    �                   �  	           `	    �                   y `	         � `	    (                   � `	          ��	    V                   Y ��	         � �"                         � po                        � 0�	    V                   	 0�	         L	  #                         p	 0p                        �	 ��	    V                   �	 ��	         
 0m     8                   C
 0�	    V                   �
 0�	         �
 �l     8                   �
 p�	    V                   ] p�	         � �#                          0q                        d ��	    V                   � ��	         4 `#                r               � �p                        � �	    V                   @ �	         � @#                         � pp     8                   D p�	    V                   � p�	         �  #                         � �o     8                    Щ	    Q                   < Щ	         p P�	    Q                   � P�	         � �	    Q                   " �	         ^ ��	    Q                   � ��	         ( Ь	    Q                   � Ь	         � �	    Q                   Y �	         � ��	    Q                   � ��	         * `    �                   k `         � �A    �                    � �A         & ��    �  	                � ��         2 P�    �  #                � P�         J  K                        �  �    7                    �         � ��    7                s         ��         � `�                      � `�         v ��    �                  � ��         f `�    F
  	                � `�         ^ `5    �  (                 `5         � p%    �  (                G p%         � H    L                  b H         � 0F    �  
                p  0F         ! ��    p                  �! ��         " P�    &                  �" P�         # ��                      �# ��          $ 0�                      �$ 0�         *% ��    �                  �% ��         4& p�    h                  �& p�         >' @�	         �' 0                         �' @                         �' �                         K(                          �( �                         �( �                         ) �                         <) p              t                 a) ��                         y) ��                        �) �                         �) �r                        �) ��                         �)  v                        �) ��                         "* ��                          M* �m                        x*  �                         �* @�     !                    �* pn                        �*  �                          +  �                          J+ ��                         n+ ��     '                    �+ �n                        �+ ��     '                    , o                        6,  �     F                    �, ��     F                    �, @�     E                    (- ��     M                    �- �n                        �- ��     !                    . 0n                        0. �[                         e. �[                     u          �. �[                         �. �[                     .text   �                       .data                           .bss    P                            �. #                         3/ T!                        p/ #                         �/ `!                        �/ #                         %0 l!                        `0 #                         �0 x!                        �0 #                         1 �!                        H1 #                         �1 �!                        �1  #                         �1 �!                        <2 $#                         w2 �!                        �2 (#                         �2 �!                        &3 ,#                         `3 �!                        �3 0#                         �3 �!                         4 4#                         34 v      �!                        f4 8#                         �4 �!                        �4 <#                         5 �!                        >5 @#                         k5 �!                        �5 D#                         �5 "                        V6 H#                         �6 "                        7 L#                         K7  "                        x7 P#                         �7 ,"                        �7 T#                         *8 8"                        |8 X#                         �8 D"                         9 \#                         q9 P"                        �9 `#                         : \"                        t: d#                         �: h"                        �: l#                         ; t"                        @; t#                         �; �"     w                         �; |#                         6< �"                        �< �#                         �< �"                        �< �#                         3= �"                        �= �#                         �= �"                        6> �#                        [> �"                        �> �#                        �> �"                        �> �#                        �> �"                        ? �#                        6? �"                        Z? �#                        �? �"                        �? �#                        �? �"                        @ �#                        :@ #                        f@ $                        �@ #                        �@ $     .                   �@ #                        2A 0B    G                     zA L$          x                      �A (#                         B T$                         DB 4#                        |B `$                         �B @#                        �B l$                         /C L#                        lC x$                         �C X#                        �C �$                         !D d#                        \D �$                         �D p#                        �D �$                         E |#                        FE �$                         �E �#                        �E �$                         �E �#                        "F �$                         SF �#                        �F �$                         �F �#                    .rdata        �  M                 �F �$     L                   G �#                        TG $%                         }G �#                 y             �G 8%                         �G �#                        �G D%                        H �#                        JH `%                        vH �#                        �H |%                        �H �#                        6I �%                        �I  $                        �I �%                        �I $                        ,J �%                        ]J $                        �J �%                         �J $$                        K �%                         <K 0$                        vK �%                         �K <$                        �K  &                         L H$                        NL &                         �L T$                        �L &                         �L `$                        6M $&                         nM l$                        z      �M (&                         �M x$                        N ,&                         KN �$                        �N 0&                        �N �$                        �N L&                        O �$                        2O h&                        |O �$                        �O �&                        P �$                        ZP �&                        �P �$                        �P �&                        �P �$                        Q �&                         XQ �$                        �Q �&                         �Q �$                        R �&                         :R �$                        nR �&                         �R �$                        �R �&                         S %                        RS '                         �S %                        �S '  {                             �S  %                        6T '                         mT ,%                        �T '                         �T 8%                        U '     (                   HU D%                        ~U D'     (                   �U P%                        �U l'     (                   KV \%                        �V �'     (                   W h%                        nW �'                         �W t%                        �W �'     (                   
X �%                        @X �'     (                   vX �%                        �X (     (                   Y �%                        nY 8(     (                   �Y �%                        0Z `(                         cZ �%                        �Z d(                         �Z �%                        :[ h(      |                         �[ �%                        �[ l(                         X\ �%                        �\ t(                         h] �%                        �] |(                         P^ �%                        �^ �(                         �^ �%                        F_ �(                         �_ &                        �_ �(                         P` &                        �` �(                         :a &                        �a �(                         b (&                        bb �(     �                   �b 4&                        �c  )     �                   d @&                        �d �)     9                   e L&                        |e �)                         f X&                        �f �)                        �f d&                        �f *             }                 �f p&                        g ,*                        [g |&                        �g H*                        �g �&                        h d*                        9h �&                        `h �*                        �h �&                        �h �*                         �h �&                        i �*                         Gi �&                        zi �*                         �i �&                        �i �*                         j �&                        .j �*                         \j �&                        �j �*     (                   �j �&                        �j �*     (                   k �&                        Jk +     (                   �k  '                         l @+     (                   [l '                        �l h+                     ~          �l '                        m l+                         �m $'                         n p+                         xn 0'                        �n t+                         Ao <'                        �o x+                         �o H'                        4p |+                         �p T'                        �p �+                         kq `'                        �q �+                         ir l'                        �r �+                         ks x'                        �s �+                         st �'                        �t �+                         wu �'                        �u �+                         Gv �'                        �v �+                         w �'                        �w �+                         )x �'                        �x �+                         ?y       �'                        �y �+                         Xz �'                        �z ,                         f{ �'                        �{ $,                         J| �'                        �| (,                         } �'                        ^} ,,                         �} �'                        N~ 0,                         �~ (                        > 4,                         � (                        � 8,                        �  (                        :� T,                        _� ,(                        �� p,                        �� 8(                        ؀ �,                        � D(                        ,� �,                         �� P(                        � �,                         R� \(                        �� �,                         � h(     �                         f� �,                         �� t(                        �� �,                        ߃ �(                        � �,                         i� �(                        ΄ �,                         	� �(                        D� �,     &                   t� �(                        �� �,     &                   ԅ �(                        � $-                         _� �(                        �� (-                         � �(                        p� ,-                        �� �(                        ʇ p�                        !� <-                          y� �(                         ш @-     &                   -� �(                        �� h-     &                   � �(                        A� �-                        e� )                        �� �-         �                     �� )                        ъ �-                         �� )                        � �-                         C� ()                        i� �-                         �� 4)                        Ջ �-                         � @)                        9� �-                         f� L)                        �� �-                        �� X)                        ی �-     (                   
� d)                        9�  .     (                   h� p)                        �� H.     (                   � |)                        K� p.     (                   �� �)                        �� �.                        +� �)                        W� �.                         �� �)                        ӏ �.                         � �)                        Q� �.                  �             �� �)                        ݐ �.                         #� �)                        i� �.                         Ց �)                        A� �.                         �� �)                        � �.                         �� �)                        � �.                         .� �)                        m� �.                         ��  *                        � �.                         � *                        [� �.                         �� *                        �  /                         J� $*                        �� /                         � 0*                        �� /                         � <*                        U� /                         �� H*                        ͘  /     <                   � T*                        Q� \/                         �      �� `*                        ٙ h/                         c� l*                        � �/                         }� x*                        � �/                         �� �*                        � �/                         �� �*                        � �/                         �� �*                        � �/                         �� �*                        � �/                         �� �*                        � 0     \                   �� �*                        [� l0     \                   � �*                        �� �0     (                   $� �*                        �� �0     4                   :� �*                        ӥ $1     h                   \� �*                        � �1     _                   n� �*                        �� �1     _                   �� +  �                            	� L2     _                   �� +                        � �2     h                   ��  +                        -� 3     h                   �� ,+                        ?� @�	    �                    �� |3                          � 8+                     .ctors  8�	                        `�  p�                          $�  ��         ��  0         �  P"         ��  0$         2�  P#         ��  �          ]�  p!         ��  �"         8�  �-         ��  )         ��  @7         @�           =� �         ��  �         �  �&         ��  �(         J�  �'         ��  %         u�  �%         	�  P'         P�  �3         �� �.         ��  0:         X�            o� �         6�  �         �           ��  �         f�           ݰ �4         }� �7         ��  P�         +�  ��        �        d�  P�         F�  ��         �  0�          ��  ��         ��  ��         )�  ��          a�  ��         ��  ��         ��  ��          �  ��         D�  p�         ~�  �          ��  p�         K�  0�         ��   �          ��  0�         ��  ��         ��  0�          �  ��         ��  �         ��  ��          �  �         ��  ��         ��  �          �  ��         ��  ��         1�  @�          i�  ��         ��  0�         �  @�          A�  0�         ��  ��         ��   �          ��  ��         �  ��         G�  `�          ��  ��         L�  ��         ��  ��          ��  ��         ��  ��         ��  ��         U�  ��         ��  ��         ��  ��          �  ��         <�  `�         �  0�         u�  @�         ��  �         ��  ��         �  `�         ;�  0�          r�  `�         V�   �         ��   �         �   �               ��   �         F�  ��         ��  `�         ��   �         ��  ��         ��               � ��    d                  �� ��         � `�    �                  �� `�         � ��                        |� ��         � �                        T� �         �� ��    �                   ;� ��         �� �    �                   1� �         �� ��    �                  5� ��         �� `�    �                  G� `�         ͹ �    K                  Y� �         ߺ `     K                  k� `          � ��    ~                   Z� ��         �� ��    ~                   &� ��         �� �                      � �         w� @�                      � @�         e� ��                        ǿ ��         #� ��                        �� ��         �� ��                    �          ]� ��         �� ��                        O� ��         �� @�    �                  v� @�         !� `�    �                  �� `�         }� ��    �                  @� ��         �� `�    �                  �� `�         }� ��    F                  /� ��         ��  �    F                  ��  �         9� Pi         $  g          \ ��          �  e          � ��           �k          @ `�          ~  k          � ��          �  i          3 ��          l  j          � ��          �  f           ��          N �g          � `�          � �e          � `�          , �l          j `�          �  l          � ��          $ �i          ] `�          � �j          � `�           �f          @ `�          �  h          � ��           �h          D `�      .text   �             �                .data                           .bss    P                            �? p�                        �? �3                          @@ D+                         �> ��                        5? �3                          x? P+                         | 0    ,                    � �3                          % \+                         z P"    n                     �3                          � h+                         J 0$    n                    � �3                          � t+                         ) P#    n                    � �3                          d �+                          �     n                    � �3                          7 �+                         � p!    n                    l  �3                          ! �+                         �! �"                        �! �3                    �            =" �+                         �" �-    �                    # �3                          �# �+                     .rdata  �     �   ,                 d�  )                       � �3     3                    �� �+                         I$ @7    n                    �$ �3                          J% �+                         �%                         & 4                          Z& �+                         �� �    #                    � 4                          �� �+                         �' �    ,                    �' 4                          I( �+                         �( �&    n                    8) 4                          �) �+                         n* �(    n                    +  4                          �+ ,                         M, �'    n                    �, (4                          �-�       ,                         &. %    n                    �. 04                          [/ ,                         �/ �%    n                    �0 84                          +1 (,                         �1 P'                        2 @4                          a2 4,                         �2 �3    �                    C3 D4                          �3 @,                         "� �.                       �� P4     3                    �� L,                         m4 0:    n                    �4 �4                          n5 X,                         �5                          66 �4                          ~6 d,                         L� �    #                    �� �4                          Y� p,                         �; �    �                    =< �4     !                    �< |,                         ��    �        �                    ]� �4     $                    �� �,                         �: �    �                    K; �4     !                    �; �,                         Y�      �                    �� 5     $                    T� �,                         �� �4                       x� (5     *                    � �,                         �� �7                       l� T5     *                    � �,                         AD P�    >                    �D �5                          �D �,                         BA ��    >                    �A �5                          �A �,                         B ��    >                    @B �5                          �B �,                         �B ��    0                    �B �5                          ?C �,                         C p�    >                    �C �5        �                         D �,                         �E 0�    >                    F �5                          FF  -                         �@ ��    0                    �@ �5                          A -                         E �    >                    CE �5                          �E -                         FG ��    <                    �G �5                          �G $-                         �F ��    <                    �F �5                          G 0-                         �I 0�    `                    �I �5                          2J <-                         xJ ��    `                    �J �5                          K H-                         �H ��    `                    I �5                          aI T-                         H ��    `                    JH �5                          �H `-               �                EN ��    F                    �N �5                          �N l-                         DQ ��    F                    �Q �5                          �Q x-                         �M ��    F                    �M  6                          N �-                         �L ��    G                    M 6                         DM �-                         IK `�    F                    �K 6                          �K �-                         R 0�    8                    ER  6                          �R �-                         L @�    F                    GL (6                          �L �-                         �P �    8                    �P 06                          Q �-                         O ��    F                    GO 86                          �O �-                         �O `�    G                  �        P @6                         FP �-                         �R  �    D                    S P6                          DS �-                         �S  �    D                    �S X6                          T �-                         U  �    h                    YU `6                          �U �-                         CT  �    h                    �T h6                          �T .                         �U ��    h                    *V p6                          pV .                         �V `�    h                    �V x6                          AW  .                         CX  �    O                    �X �6                         �X ,.                         �W ��    O                    �W �6                         X 8.                         �� �6     <                   :� D.                        �� �6�           L                   :� P.                        �� (7                         *� \.                        �� ,7                         
� h.                        z� 07     !                   �� t.                        x� T7     !                   �� �.                        v� x7     G                   � �.                        �� �7     G                   � �.                        �� 8     ]                   7� �.                        �� h8     ]                   Q� �.                        �� �8                         H� �.                        �� �8                         � �.                        �� 9     +                   � �.                        |� 49     +                   �� �.                        r� `9                         �� �.                        8� d9     �                          �� �.                        �� h9                         {� /                        �� l9                         u� /                        �� p9                         �� /                        V� x9                         � (/                        �� �9     ,                   ~� 4/                        B� �9     ,                   � @/                        �� �9     /                   }� L/                        0� :     /                   �� X/                        �� Pi    ;	  q                 �� 8:     �                    �� d/                         ww  g     8                    �w ��     5                     �w  e     8                    3x ��     4                     qx �k     8                    �x `�     ;                     �x  k     8                    @y ��     ;       �                    �y  i     8                    �y ��     6                     z  j     8                    Ez ��     6                     �z  f     8                    �z ��     5                     { �g     8                    B{ `�     5                     �{ �e     8                    �{ `�     4                     �{ �l     8                    B| `�     ;                     �|  l     8                    �| ��     ;                     } �i     8                    Q} `�     6                     �} �j     8                    �} `�     6                     ~ �f     8                    P~ `�     5                     �~  h     8                    �~ ��     5                      �h     8                    L `�     5                     � @�     H                    � 0�     8                    � `�     h                    M� ��     h              �            �� ��     0                    Ҁ ��     0                    � 0�     8                    Q� �     H                    �� ��     8                    ΁  �     h                    � @�     h                    X�  �     0                    �� �     0                    ؂ ��     8                    � ��     X   
                 V� 0�     X   
                 +� p    	                    g� p                          ��  �    	                    ��  �         � `                        I� `         }� �}                        �� �}         �� �}                        "� �}         U� ��    	                    �� ��         �� `�    	                    � `�         9� ��                        s� ��         �� 0�                        �� 0�         �  �                        L�  �         � P-	        �                     �� P-	         ��  �     h                   �  1	                       A�  1	         m� p�     h                   ��  �    	                    ��  �         � 0�    	                    8� 0�         g� @ 	                       �� @ 	         �� �     H                   �� 0�                        C� 0�         �� �                        �� �         [�  �                        ��  �         �� `�    "                    �� `�         � `A	                       V� `A	         �� p�     0                   �� �B	                       C� �B	         �� ��     0                   �� @@	                       /� @@	         y� �     X   
                �� �!	                       !  �!	         s   -	    $                   �   -	         �  �0	    $                    �0	         / 0A	  �        $                   � 0A	         � PB	    $                    PB	         g  	    $                   �  	         � @	    $                   	 @	         S �!	    $                   � �!	         � �7	    (                   ! �7	         ? ��     8                   c �7	    0                   � �7	         � @4	    (                   � @4	         �  �     8                    4	    0                   + 4	         H `	    (                   t `	         � 0	    0                   � 0	         � @	    (                    @	         < 	    0                   g 	         � ��    &  	                � ��         � �C         : p�    H                   q p�         � 0}    H                   � 0}         
 Э    H                   : Э         d ��    H   �                      � ��         � P�    H                   	 P�         D	 �    H                   �	 �         �	 p�    H                   �	 p�         
     H                   L
          �
  �    H                   �
  �         �
 �    H                    �         L �    H                   � �         � �    :                  � �         ��              " �    L                   M �         r �     h                   �  �    L                   �  �         � P�    H                   6 P�         y `�    H                   � `�          ��    G                   5 ��         _ ��    G                   � ��         � �}    #                   � �}         % �~    #                   ^ �~         � 0�    o                   � 0�         � �| �         o                   ( �|         Y p~    o                   � p~         �  ~    o                   �  ~         1 �}    #                   h �}         � �|    #                   � �|         � `|    #                   5 `|         e ��    L                   � ��         � P�     h                   � и    L                    и         0  �    H                   y  �         � 0�    H                    0�         H p�    G                   x p�         � ��    G                   � ��         � ��    #                   5 ��         h  �    #                   �  �         � p�    o                    p�         4  �    o                   k  �         � ��    o                   � ��          @�    o                   A @�         t ��    # �                        � ��         � Ѐ    #                    Ѐ         B ��    #                   x ��         � `+	    �                   � `+	          �)	    �                   A �)	         p @,	    �                   � @,	         * �*	    �                   � �*	         � `-	                        `-	         B 0/	    �                   w 0/	         � p-	    �                   � p-	         
 0	    �                   j 0	         � P.	    �                   $ P.	         ~ 01	                       � 01	         � A	                       - A	         x �@	                       � �@	          0i    k                    � 0i            �h    k                    �  �h         $! pA	                       u! pA	         �! 0B	                       " 0B	         \" B�      	                       �" B	         �" ��    ^                    ]# ��         �#  �    S                    ?$  �         �$ �B	                       % �B	         X% ��    �  -                �% ��         t& �"                         �&  �    �  -                0'  �         �' �"                         �' @�    �                  N( @�         �( ��    ^                   6) ��         �) p>	    I                   �) p>	         �) 0�     H                   * �=	    I                   @* �=	         ^* �=	    E                   �* �=	         �* �<	    E                   + �<	         B+  >	    G                   h+  >	         �+ 0=	    G                   �+ 0=	         �+ ��    #                    , ��         ,, �    #                   ^, �         �, @�    o                   �, @�     �          �, ��    o                   - ��         .-  �    o                   [-  �         �- P	    �                   �- P	         �- �	    �                   	. �	         2. 0	    �                   �. 0	         �. p	    �                   :/ p	         �/ P 	                       �/ P 	         �/ �6                       Z0 �6         �0 �Q                        $1 06                       �1 06         2 �?	                       b2 �?	         �2 �?	                       �2 �?	         F3 ��    #                   �3 ��         �3 �$    _                    t4 �$         �4 P$    _                    j5 P$         �5 ��    _                    d6 ��         �6 @�    _                    d7 @�         �7 %    _                    `8 %         �8 P@	                       (9 P@	         r9 �      ��    �                  �9 ��         x: ��    �                  �: ��         v; �    �                  < �         �< ��    �                  = ��         �= �    K                  > �         �> p!	                       �> p!	         P? ��     X   
                �? 0!	                       @ 0!	         X@ �!	                       �@ �!	         FA P!	                       �A P!	         4B �!	                       �B �!	         �B `7	    B                   C `7	          C �6	    B                   DC �6	         bC 7	    B                   �C 7	         �C p6	    B                   �C p6	         �C @�    #                   ZD @�         �D p�    #                   E p�         tE �    ,                    �E �         F ��                       EF ��         hF 8	    �      (                   �F 8	         �F �                        G �         lG �                        �G �         �G p	    �   
                	H p	         2H ��     8                   ^H �	    �   
                �H �	         �H  	                       I  	         dI `	                       �I `	         J �	    (                   >J �	         dJ ��         �J ��         K @	    �                   aK @	         �K 0Q                        �K `    �                   <L `         �L �3	    B                   �L �3	         �L 03	    B                   �L 03	         M �3	    6                   6M �3	         UM �2	    6                   zM �2	         �M P�                        �M P�         �M ��                        .N ��         YN  �    #                   �N  �         �N�       p4	    (                   �N p4	         �N P	    �                   O P	         AO  �     8                   lO �	    �                   �O �	         �O 0	    �                   P 0	         nP p	    �                   �P p	         Q p	    (                   EQ p	         jQ �	    V                   �Q �	         �Q �"                         R �o                        $R ��	    V                   bR ��	         �R 0#                         �R Pp                        �R P�	    V                   'S P�	         fS �m     8                   �S �	    V                   �S �	         T pm     8                   @T н	    V                   �T н	         U �#                         aU Pq                        �U �	    V                   V �	         �V p#                         �V q   �                           $W P�	    V                   �W P�	         �W P#                         BX �p     8                   �X к	    V                   �X к	         Y #                         ,Y �o     8                   PY 0�	    Q                   �Y 0�	         �Y ��	    Q                   �Y ��	         .Z p�	    Q                   pZ p�	         �Z �	    Q                   [ �	         v[ 0�	    Q                   �[ 0�	         @\ p�	    Q                   �\ p�	         ] �	    Q                   C] �	         x] `    �                   �] `         �] �B    �                    7^ �B         t^ @�    �                  �^ @�         �_ `�    �                  ` `�         �` 0K                        �` `�    �                  Ta `�         �a ��    �                  Rb ��         �      �b P"    �                  Lc P"         �c �    �                  ?d �         �d Y    �  '                \e Y         �e `I    �  '                �f `I         Hg pk    {                  �g pk         :h �i    �                  �h �i         di 0H    
                  �i 0H         nj �a    r  
                �j �a         xk P;    �  
                 l P;         �l @U    `  
                
m @U         �m  n    >  
                n  n         �n `{    �  
                o `{         �o �    �                  p �         �p ��	         �p P                         %q `                         Rq                           �q                           �q �                         r �                         pr �                         �r �                         �r ��  �                             �r ��                          	s n                        4s  �                         Xs ��     !                    �s �n                        �s `�                          �s @�                          t ��                         *t  �     '                    \t 0o                        �t @�     '                    �t Po                        �t `�     F                    Cu  �     F                    �u ��     E                    �u  �     M                    <v �n                        �v  �     !                    �v Pn                        �v \                         !w  \                         Vw �[                         �w �[                     .text   �                       .data                           .bss    P                            �w �:                         �w p/      �                        ,x �:                         ix |/                        �x �:                         �x �/                        y �:                         Vy �/                        �y �:                         �y �/                        z  ;                         Az �/                        ~z ;                         �z �/                        �z ;                         3{ �/                        n{ ;                         �{ �/                        �{ ;                         | �/                        V| ;                         �| �/                        �| ;                         �| �/                        "} ;                         X}  0                        �}  ;                         �} 0                        �} $;                         '~ 0             �                 T~ (;                         �~ $0                         ,;                         v 00                        � 0;                         � <0                        4� 4;                         d� H0                        �� 8;                         � T0                        8� <;                         �� `0                        ܁ @;                         -� l0                        ~� D;                         ׂ x0                        0� H;                         c� �0                        �� P;                         Ƀ �0                        �� X;                         N� �0                        �� `;                         � �0                        D� h;                         q� �0                        �� p;                         � �0                    �          @� x;                         �� �0                        � �;                        � �0                        <� �;                        a� �0                        �� �;                        �� �0                        · �;                        � �0                        � �;                        C� 1                        p� �;                        �� 1                        ʈ �;                        ��  1                        "� �;                        N� ,1                        z�  <     .                   �� 81                        � �C    H                     6� 0<                          � D1                         Ȋ 8<                          � P1                        8� D<                         p� \1                        �� P<                         ً �      h1                        
� \<                         G� t1                        �� h<                         �� �1                        �� t<                         7� �1                        t� �<                         �� �1                        ؍ �<                         � �1                        N� �<                         � �1                        �� �<                         � �1                        *� �<                         g� �1                    .rdata  �	     �  M                 �� �<     X                   ڏ �1                        � =                        <� �1                        h� 0=                        �� �1                        �� L=                        
� �1                        T� h=                        �� 2                        � �=     �                         � 2                        J� �=                        {� 2                        �� �=                         � (2                         � �=                         Z� 42                        �� �=                         ȓ @2                        �� �=                         4� L2                        l� �=                         �� X2                        �� �=                         � d2                        T� �=                         �� p2                        ĕ �=                         �� |2                        2� �=                         i� �2                        ��  >                        ̖ �2                        �� >                        $� �2                        P� 8>                        �� �2                        � T>         �                     .� �2                        x� p>                        �� �2                        ژ �>                        � �2                        <� �>                         v� �2                        �� �>                         � �2                        $� �>                         X� �2                        �� �>                         Ě  3                        �� �>                         6� 3                        p� �>                         �� 3                        � �>                         � $3                        T� �>                         �� 03                         �>                         �� <3                        0� �>     (                   f� H3                        �� ?     (                   ҝ T3                        � <?     (            �             i� `3                        ʞ d?     (                   +� l3                        �� �?                         �� x3                        � �?     (                   (� �3                        ^� �?     (                   �� �3                        ʠ �?     (                   +� �3                        �� @     (                   � �3                        N� 0@                         �� �3                        �� 4@                         � �3                        X� 8@                         �� �3                        �� <@                         v� �3                        � D@                         �� �3                        � L@                         n� �3                        �� P@                         � �3                        d� T@                         �      �� 4                        � X@                         n� 4                        Ԩ `@                         X�  4                        ܩ h@                         .� ,4                        �� l@     �                   � 84                        �� �@     �                   6� D4                        Ȭ �A     9                   1� P4                        �� �A                         !� \4                        �� �A                        ͮ h4                        � �A                        � t4                        <� B                        y� �4                        �� $B                        � �4                        0� @B                        W� �4                        ~� \B                        �� �4                        ̰ xB                         �� �4  �                            2� |B                         e� �4                        �� �B                         ű �4                        � �B                         � �4                        L� �B                         z� �4                        �� �B     (                   ز �4                        � �B     (                   8� �4                        h� �B     (                   ó 5                        � C     (                   y� 5                        Դ DC                         � 5                        .� HC                         �� (5                        $� LC                         �� 45                        � PC                         k� @5                        �� TC                         � L5                        ^� XC                         �� X5      �                        � \C                         �� d5                        � dC                         �� p5                        � lC                         �� |5                        � tC                         �� �5                        "� |C                         �� �5                         � �C                         q� �5                        ¾ �C                         I� �5                        п �C                         S� �5                        �� �C                         i� �5                        �� �C                         �� �5                        � �C                         �� �5                        �  D                         t� �5                        �� D                         ,� �5                        �� D                         �  6             �                 ~� D                         �� 6                        t� D                         �� 6                        &� D                        K� $6                        p� 0D                        �� 06                        �� LD                        �� <6                        � hD                        8� H6                        b� �D                         �� T6                        $� �D                         �� `6                        �� �D                         D� l6                        �� �D                         �� x6                        �� �D                        � �6                        :� �D                         �� �6                        � �D                         ?� �6                        z� �D     &                   �� �6                    �          �� �D     &                   
� �6                        :�  E                         �� �6                        �� E                         K� �6                        �� E                        �� �6                         � ��                        W� E                          �� �6                         � E     &                   c� �6                        �� DE     &                   � �6                        w� lE                        �� 7                        �� �E                        �� 7                        � �E                         -�  7                        S� �E                         y� ,7                        �� �E                         �� 87                        � �E                         =� D7                        o� �E                         �� �      P7                        �� �E                        �� \7                        � �E     (                   @� h7                        o� �E     (                   �� t7                        �� $F     (                   '� �7                        �� LF     (                   �� �7                        5� tF                        a� �7                        �� �F                         �� �7                        	� �F                         H� �7                        �� �F                         �� �7                        � �F                         Y� �7                        �� �F                         � �7                        w� �F                         �� �7                        O� �F                         �� �7                        %� �F                         d� �7     �                         �� �F                         �� 8                        � �F                         U� 8                        �� �F                         �� 8                        � �F                         �� (8                        �� �F                         R� 48                        �� �F                         #� @8                        �� �F                         �� L8                        � �F     <                   E� X8                        �� 8G                         �� d8                        � DG                         �� p8                        #� \G                         �� |8                        C� tG                         �� �8                        I� �G                         �� �8                        O� �G                         �� �8         �                     M� �G                         �� �8                        E� �G     `                   �� �8                        �� 8H     `                   @� �8                        �� �H     (                   f� �8                        �� �H     4                   |� �8                        � �H     T                   �� �8                        '� HI     S                   �� �8                        9� �I     S                   ��  9                        K� �I     S                   �� 9                        ]� DJ     S                   �� 9                        o� �J     S                   �� $9                        �� �J                         � 09                        �� ��	    �                    �� K                          ^� <9                     .ctors  @�	                �              �� ��                       � ��                          I� `�    ,                   �� `�         �� `�                       � `�         A� 0�    ,                   �� 0�         �� ��                       � ��         A� ��    !                   �� ��         �� ��    4                   � ��         Y� ��    	                   �� ��         �� ��    	                   � ��         ]� P�    7                   �� P�         �� P�    m                   O� P�         �� ��    m                   � ��         {� ��                       �� ��         �� �    u                   G� �         �� `�    "                   �� `�         �  �    7                   ^�  �         �� ��    7                   �� ��         +� ��    I                   t� ��         �� 0�       �                         0�         C  ��    6                   �  ��         �  P�    �                   . P�         � ��    �                   � ��         E ��    @                   � ��         � �P                        � ��    @                   - ��         c �P                        � ��    H                   � ��          ��    H                   K ��         � `�                       � `�         � 0�     �                   / �                       k �         � ��    �                   � ��         7 0�    �                   � 0�         �  �    �                   "  �         q ��    �                   � ��          �    @                   Q �         � p�                       � p�         	 P�    	                   B	 P�         y	 `� �         	                   �	 `�         �	 ��    o                   9
 ��         {
 0�     �                   �
 @�    o                    @�         F ��    ?                   � ��         �  �    ?                     �         J ��    8                   � ��         � ��    �                    ��         T ��                        � ��         � `�                        `�         H ��     �                   � ��                       � ��         � ��    �                   D ��         � 0�    �                   � 0�         "  �    �                   w  �         � ��    �                    ��         j �    @                   � �         � p�                        p�         Z P�    	                   � P�         � `�    	                 �         `�         F ��    q                   � ��         � ��     �                    ��    q                   Y ��         � `�    C                   � `�          ��    C                   a ��         � ��    <                   � ��         !  �    �                   h  �         � ��                        � ��         +  �     6                    l  d                        � `�     6                    �  d                        / ��     1                    k �c                        � ��     1                    � �c                    .text   �                       .data                           .bss    P                             K                         a H9                        � K                         � T9                        ' K                         i `9�                              � K                         � l9                        /  K                         u x9                        � (K                          �9                        O 0K                         � �9                        � 8K                         ( �9                        m <K                         � �9                        � @K                         @ �9                        � HK                         � �9                        [ TK                         � �9                        -  `K                         s  �9                        �  hK                         ! �9                        K! xK                         �! �9                        �! �K                         )" �9                        s" �K                         �" :     �                         # �K                         O# :                        �# �K                         �#  :                        -$ �K                         v$ ,:                        �$ �K                         !% 8:                        �% �K                         �% D:                        G& �K                        �& P:                        �& �K                        �& \:                        ;' �K                        x' h:                        �' �K                        �' t:                        /( L                         l( �:                        �( L                         �( �:                        #) L     &                   r) �:                        �) @L     &                   * �:                        _* hL     &                   �* �:           �                   + �L     &                   a+ �:                        �+ �L                        �+ �:                        1, �L                         t, �:                        �, �L                         �, �:                        3- �L                         s- �:                        �- �L                         �- �:                        E. �L                         �. ;                        �. �L                        / ;                        a/  M                        �/ ;                        �/ M                        00 (;                        u0 (M                         �0 4;                        1 8M                         J1 @;                        �1 <M                         �1 L;                        	2 DM                         F2 X;                  �            �2 LM     &                   �2 d;                        !3 tM     &                   p3 p;                        �3 �M     &                   4 |;                        k4 �M     &                   �4 �;                        5 �M                        T5 �;                        �5 �M                         �5 �;                        6  N                         U6 �;                        �6 N                         �6 �;                        7 N                         \7 �;                        �7 N                         �7 �;                        78  N                        |8 �;                        �8 4N                        9 �;                        K9 HN                        �9 �;                        �9 \N                         :  <                        e:�       lN                         �: <                        �: �    ]                   *; �                          _; 7    ]                   �; 7         �; �    �                   < �         A< PA    �                   }< PA         �< `    +                    �< `         = �3    ,                    R= �3         �= p0         �= �    .                   > �         F>  @    A                   �>  @         �> �    0                  �> �         *?  B                      f?  B         �? P    .                  �? P         @ �9    >                  J@ �9         �@     3                  �@          �@ p7                      +A p7         `A �	    ;                    �A �	         �A �	    D                    $B �	         bB @(    N  	                �B @(  �             �B �     �                   �B P%    N  	                *C P%         XC �&    �                  �C �&         �C �#    �                  �C �#         (D P                      bD P         �D �:    	                   �D �:         E      3                   UE           �E �    k                   �E �         4F      e                  �F           �F  	    r                    	G  	         FG 
                      �G 
         �G �    �                   H �         ^H �    �                  �H �         �H @    �                  )I @         ~I     �                   �I           J �                      bJ �         �J �    k                    �J �         K ��                      RK ��         �K ��    S  	                �K ��         �      �K  a     P                   %L ��     P                   XL ��    �                   �L ��         �L P;                        M P;         6M ��    	                   qM ��         �M `;    	                   �M `;         N ��    �                   PN ��         �N �    ;  	                �N �         �N @b     P                   #O  �     P                   VO �    �                   �O �         �O �;                         P �;         4P  �    	                   oP  �         �P �;    	                   �P �;         Q �V    m                  MQ �V         ~Q  Q    f  
                �Q  Q         �Q @_     P                   R �     x   	                NR �_     P                   �R P    �                   �R P         �R �:                        ,S �:         _S Q �         	                   �S Q         �S �:    	                   T �:         =T �,    ;                    �T �,         �T -    G                    U -         ?U �K    S  	                sU �K         �U ��     �                   �U �H    S  	                V �H         5V  J    �                  lV  J         �V  G    �                  �V  G         W �1                      ?W �1         sW �:    	                   �W �:         �W P0                       2X P0         {X �/    k                   �X �/         Y p.    e                  ]Y p.         �Y P,    u                    �Y P,         #Z `-                      jZ `-         �Z �:    �                   �Z �:         ;[  >    �                  v[  >         �[ �;    �                  \ �;         [\ P=    � �                        �\ P=         �\ �4                      ?] �4         {] �+    k                    �] �+         �] ��                      /^ ��         a^ ��    [  	                �^ ��         �^ Pa     P                   _ 0�     P                   J_ `�    �                   �_ `�         �_ p;                        �_ p;         (` p�    	                   c` p�         �` �;    	                   �` �;         
a �    �                   Ba �         ta  �    C  	                �a  �         �a �b     P                   *b P�     P                   ]b �    �                   �b �         �b �;                        c �;         ;c �    	                   vc �         �c �;    	                   �c �;         d �f    n                  Td �f         �d �`    n  
     �                 �d �`         �d �_     P                   8e ��     x   	                je �`     P                   �e �_    �                   �e �_         $f �:                        ]f �:         �f �`    	                   �f �`         �f  ;    	                   9g  ;         ng ��	    ^                   �g ��	         h �    �                   >h �         ph  *    <                   �h  *         �h �)    <                   i �)         4i ��    �                   ii ��         �i ��       
                �i ��         �i ��    �                   1j ��         `j ��    �   
                �j ��         �j  [                      �j  [         &k �U    3                  Zk �U         �k `*                      �k `*         �k ��    �                   (l ��         Zl @^    �      �                   �l @^         �l ��    �                   �l ��         ,m @    �                   vm @         �m @                       (n @         �n P�    J                   �n P�         ho ��    J                   �o ��         @p �O    G                   �p �O         q  �    G                   aq  �         �q p�    G                   �q p�         6r pO    G                   �r pO         �r �R    �                  s �R         Ls `X    ]  	                �s `X         �s  T    �                  ?t  T         �t �Y    ^  	                u �Y         tu ��    �                   �u ��         �u ��    �                   Fv ��         �v �    N                  �v �         w P�    8                  Zw P�         �w ��    �                   x ��         nx �      ��    �                   �x ��         @y ��    C                  �y ��         z `�    N                  ~z `�         �z `�    :                   { `�         P{ ��    :                   �{ ��         �{ �P    :                   �{ �P         &| p�    u                   [| p�         �| @�    m                   �| @�         �| ��       	                #} ��         R} ��    �   	                �} ��         �} �\    �   
                �} �\         ~ �)    D                   L~ �)         z~  �	    �   	                �~  �	         �~ 0�	    �   	                + 0�	         b ��	    �   
                � ��	         � ��	    �   
                � ��	         B� �]    �                   v� �]         �� @\    �                   ؀ @\         � P�    �   
                ;� P�    �           j� 0�    �   
                �� 0�         ΁ ��	    �   
                � ��	         B�  �	    �                   |�  �	         �� ��	    �   
                � ��	         $� ��	    �                   `� ��	         �� 0�	    ^                   � 0�	         .� �3    �                   f� �3         �� �M    <                   ̄ �M         �� pM    <                   .� pM         \� ��    �                   �� ��         �� ��      
                �� ��         $� ��    �                   Y� ��         �� �    �   
                �� �         � �j                       � �j         N� `e    :                  �� `e         �� �M                      � �M         � ��    �                   P� ��         �� �m    �                   �� �m         � �    �                   "��       �         T� �0    �                   �� �0         � �1                       S� �1         �� �    J                   0� �         �� ��    J                   � ��         z� `_    G                   � `_         V� ��    G                   �� ��         � p�    G                   1� p�         v� _    G                   �� _         � @b    �                  K� @b         �� h    ]  	                ӏ h         � �c    �                  �� �c         � pi    ^  	                X� pi         ��  �    �                   �  �         J� ��    �                   �� ��         Ԓ p�    C                  � p�         ^� ��    R                  �� ��         � ��    �                   W� ��         �� ��    �                   /� ��         �� ��    C           �             � ��         p� @�    S                  ߖ @�         H� 0�    :                   �� 0�         �� ��    :                   � ��          � �`    :                   X� �`         �� �    m                   �� �         � p�    u                   #� p�         R�         	                ��           �� ��    �   	                � ��         � �l    �   
                N� �l         |�  M    D                   ��  M         ޚ ��	    �   
                � ��	         P� @�	    �   	                �� @�	         ě  �	    �   
                ��  �	         2� `�	    �   	                o� `�	         �� @m    �                   ڜ @m         � �k    �                   <� �k         j� p     �   
                �� p          Ν P�    �   
                � P�         2� ��	    �   �      
                o� ��	         �� @�	    �                   � @�	         � ��	    �   
                U� ��	         �� p�	    �                   Ɵ p�	         �� ��                          %� �b                        P�  �     '                    ��  u                        �� ��     (                    � 0v                        � ��     (                    M� �v                        �� ��     '                    �� `u                        � `�     '                    � @u                        H�  �     (                    {� Pv                        �� ��     (                    � �v                        � ��     '                    F� �u                        x�  �                         �� ��                         ޣ �^     x                   � @�     P   
                F�  �                �               y� ��                         �� 0`     x                   �� ��     P   
            .text   �                       .data                           .bss    P                            *� pN                         f� <                        �� |N                         ޥ $<                        � �N                         W� 0<                        �� �N                         Ѧ <<                        � �N                         F� H<                        ~� �N                         �� T<                        � p0    7                    E� �N                          �� `<                         �� �N                         2� l<                        o� �N                         �� x<                    .rdata  �     G                    � �N                         &� �<                      �        c� �N                         �� �<                        ݪ  O                         � �<                        W� O                         �� �<                        ѫ  O                         � �<                        I� 0O                         �� �<                        �� @O                         � �<                        I� DO                         �� �<                        ӭ HO     #                   � �<                        =� lO     #                   r� �<                        �� �O                         ߮ �<                        � �O                         O� =                        �� �O                         ¯ =                        �� �O                         9�  =                        u� �O                         Ű ,=                        � �O�                               d� 8=                        �� �O                          � D=                        M� �O                         �� P=                        ղ �O                         � \=                        e� P                         �� h=                        �� P                         9� t=                        u� $P                         Ѵ �=                        -� 8P                         �� �=                        ׵ HP                         � �=                        ]� TP                         �� �=                        � XP     '                   � �=                        S� �P     )                   �� �=                        ŷ �P                        � �=                        =� �P                         x� �=                        �� �P     �                          � �=                        +� �P                         h� �=                        �� �P     '                   ޹ �=                        � �P     )                   P� >                        �� $Q                        ź >                        � <Q                         <� >                        w� @Q                         �� (>                        � DQ                         ,� 4>                        i� HQ     '                   �� @>                        ټ pQ     )                   � L>                        I� �Q                        �� X>                        �� �Q                         �� d>                        3� �Q                         n� p>                        �� �Q                         � |>                        !� �Q            �                   e� �>                        �� �Q                         � �>                        3� �Q     #                   h� �>                        �� �Q     #                   �� �>                        � R                         ?� �>                        w� R                         �� �>                        �� (R                         "� �>                        ]� 8R                         �� �>                        �� <R                         %� �>                        u� @R                         �� �>                        � HR                         `�  ?                        �� `R                         �� ?                        5� lR                         }� ?                        �� �R                         � $?                        ]� �R                   �            �� 0?                        �� �R                         1� <?                        �� �R                         �� H?                        7� �R                         z� T?                        �� �R                         �� `?                        A� �R     '                   z� l?                        �� �R     )                   �� x?                        %� (S                        a� �?                        �� @S                         �� �?                        � DS                         O� �?                        �� HS                         �� �?                        � LS     '                   >� �?                        w� tS     )                   �� �?                        �� �S                        %� �?                        a� �S                         ���       �?                        �� �S                         � �?                        O� �S                         �� �?                        �� �S     '                   � �?                        9� �S     )                   q� @                        �� T                        �� @                        � 0T                         Y�  @                        �� 4T                         �� ,@                        	� 8T                         E� 8@                        �� <T                         �� D@                        !� DT     <                   Z� P@                        �� �T                        �� \@                        �� �T                        2� h@                        g� �T     *                   �� t@                        �� �T     .                   	� �@   �                           ?� �T     (                   u� �@                        �� $U     .                   �� �@                        � TU     2                   L� �@                        �� �U     9                   �� �@                        �� �U                         #� �@                        [� �U                        �� �@                        �� �U                        � �@                        =� V                        v� �@                        �� 0V                         �� �@                        E� @V                         �� �@                        #� DV                         �� A                        � LV                         s� A                        �� TV                         R� A                        �� \V                         � (A        �                      Y� dV                         �� 4A                        �� lV                         <� @A                        �� tV     9                   �� LA                        � �V     2                   _� XA                        �� �V     9                   � dA                        �  W     2                   �� pA                        W� TW     +                   �� |A                        �� �W     +                   2� �A                        {� �W     3                   �� �A                        � �W     2                   V� �A                        �� X     +                   � �A                        y� @X     +                   �� �A                        S� lX     2                   �� �A                        -� �X     3                   �� �A               �               � �X                         A� �A                        {� �X                         �� �A                        �� �X                         (� �A                        a� �X                        ��  B                        ��  Y                        � B                        9� Y                        o� B                        �� $Y                        �� $B                        � 4Y                        F� 0B                        {� DY                        �� <B                        �� TY                        #� HB                        a� dY                        �� TB                        �� tY                        � `B                        W� �Y                        �� lB                        �� �Y                        � xB                      �        7� �Y                        l� �B                        �� �Y                        �� �B                        � �Y                        C� �B                        y� �Y                        �� �B                        �� �Y                        0� �B                        k� �Y                        �� �B                        �� Z                        $� �B                        a� Z                         �� �B                        � $Z     <                   :� �B                        s� `Z                        �� �B                        �� pZ                        � �B                        G� �Z     *                   }� C                        �� �Z     /                   �� C                        � �Z     (                   U�  C                        �� [�           .                   �� ,C                        �� 4[     2                   ,� 8C                        a� h[     9                   �� DC                        �� �[                         � PC                        ;� �[                        t� \C                        �� �[                        �� hC                        � �[                        V� tC                        �� \                         �� �C                        %�  \                         �� �C                        	� $\                         |� �C                        �� ,\                         b� �C                        �� 4\                         G� �C                        �� <\                         � �C                        Q� D\                         �� �C                        �� L\     �                          4� �C                        � T\     9                   �� �C                        � �\     2                   W� �C                        �� �\     9                   � �C                        }�  ]     2                   �� D                        [� 4]     +                   �� D                        �� `]     +                   6� D                        � �]     3                   �� (D                          �]     3                   Z  4D                        �  �]     +                    @D                        �  ^     +                   � LD                        c L^     3                   � XD                        C �^     3                   � dD                        # �^                         ] pD                        � �^            �                   � |D                         �^                         D �D                        } �^                        � �D                        � �^                         �D                        U �^                        � �D                        � _                        � �D                        - _                        b �D                        � $_                        � �D                         4_                        > �D                        { D_                        � �D                        � T_                        2	 �D                        m	 d_                        �	  E                        �	 t_                        
 E                        S
 �_                        �
 E                        �
 �_                  �            �
 $E                        ) �_                        _ 0E                        � �_                        � <E                         �_                        N HE                        � �_                        � TE                         �_                        B `E                        } `                         � Т	                          � �P                        �  u                        � ��	          pS                        # ��                        ; @�	         S  S                        r                          � P�	         �  P                        � Pr                        �  �	         � �s                         ��	         5 `t                        Q �	         s y                        � 0�	         � �t         �                     � ��	         � �t                         `�	         * �	         I v                        f p�	         � �s                        � `�	         � pw                        � ��	         � �x                          �                         9 ��                         P �                         j  �                         � ��                         � `�                         � ��                         � ��                         � ��                          ��                         . �                         I ��                         g @�                         �  K                        � �J                        � �J                        � �J                        ' �J                        N �J                        u K                 �             � �J                        � �J                        � �I                         `M                        4 N                        W �J                    .text   �                       .data                           .bss    P                             Т	    3                    � �_                          � lE                         � ��	    3                    	 `                          ) xE                         I @�	    3                    g `                          � �E                         � P�	    3                    � `                          � �E                           �	    K                    * `                         N �E                         r ��	    K                    � 8`                         � �E                         � �	    K                    �       T`                         1 �E                         Z 0�	    K                    ~ p`                         � �E                         � ��	    K                    � �`                          �E                         6 `�	    �   
                 _ �`     $                    � �E                         � �	    K                    � �`                         � �E                         $ p�	    K                    G �`                         k �E                         � `�	    K                    � a                         � �E                          ��	    K                    *  a                         R F                         L�                               ��              z @|	                       � @|	         �  �                         �  �	                       .  �	 �              W  �                         � |	    $                   � |	         � ��	    $                    ��	         4 ��                        e ��         � Є                        � Є         � ��                          ��         P Pv	    2                   � Pv	         � z	                        z	         R  s	                       �  s	         � ��    	                     ��         > ��    	                    p ��         �  �                        �  �         � Ђ                        .  Ђ         Z  ��                        �  ��         �  s	                       ! s	         R! P|	                       �! P|	         �! ��                        �! ��         " �s	                        ;" �s	         h" ��                        �" ��       �        �" @w	    5                   # @w	         \# �    �                   �# �         �# �s	    �                   �# �s	         $ 0�    l                   P$ 0�         �$ ��    c                   �$ ��         �$ �{	    ]                   % �{	         :% �z	    ]                   i% �z	         �%  z	                        �%  z	         ,& @s	    �                   t& @s	         �& �w	    �                  �& �w	         "' �v	    �   
                _' �v	         �' �t	    T                   �' �t	         &(  {	    �                   n(  {	         �( 0z	    �                   �( 0z	         :) Pu	    e                   o) Pu	         �) �u	    �                   �) �u	         * �t	    e                   7* �t	         f* 0�                        �* 0�         �* @�                        �* @��               + �                        R+ �         �+ p	    2                   �+ p	          , Ђ	                       E, Ђ	         �, p|	                       �, p|	         - ��    	                    C- ��         p-  �    	                    �-  �         �-  �                        .  �         .. ��                        `. ��         �. ��                        �. ��         �. `|	                       B/ `|	         �/ 0�	                       �/ 0�	         �/ �                        0 �         :0  }	                        �0  }	         �0 ��                        �0 ��         &1 `�	    5                   r1 `�	         �1 0�    Q                   �1 0�         2 0}	    b                   J2 0}	         v2 ��    +                   �2 ��         �2 ��    '               �          3 ��         >3 ��	    d                   m3 ��	         �3 ��	    d                   �3 ��	         �3 ��	                        >4 ��	         �4 �|	    �                   �4 �|	         5 ��	    $                  K5 ��	         ~5 �	    �   
                �5 �	         �5 �}	    [                   =6 �}	         �6 ��	    �                   �6 ��	         7 ��	    �                   T7 ��	         �7 p~	    f                   �7 p~	         �7 �~	    �                   /8 �~	         ^8  ~	    f                   �8  ~	         �8 ��                         �8                          �8  �     "                    9 Ѐ                        J9 `�     "                    w9 ��                    .text   �                       .data                           .bss    P                            �9 <a            �                   �9 F                        : @a                         4:  F                        d: Da                         �: ,F                        �: La                         �: 8F                        $; Ta                         V; DF                        �; Xa                         �; PF                        �; \a                         !< \F                    .rdata  �                          X< `a                         �< hF                        �< ha                         $= tF                        j= la                         �= �F                        �= ta                         2> �F                        f> xa                         �> �F                        �> |a                          ? �F                        4? �a                         g? �F                  �            �? �a                         �? �F                        @ �a                         Y@ �F                        �@ �a                         �@ �F                        A �a                         5A �F                        hA �a                         �A �F                        �A �a                         B �F                        :B �a                         �B G                        �B �a                         C G                        <C �a                         oC G                        �C �a                         �C (G                        D �a                         ED 4G                        zD �a                         �D @G                        �D �a                         
E LG                        :E �a                         �E XG                        �E�       �a                         %F dG                        nF �a                         �F pG                        �F b     '                    G |G                        ^G ,b                         �G �G                        �G 8b                        ?H �G                        �H Tb                        �H �G                        I pb                         PI �G                        �I |b                        �I �G                        �I �b                         (J �G                        ^J �b                         �J �G                        �J �b                         �J �G                        $K �b                         [K �G                        �K �b                         �K �G                        L �b                         ^L  H                        �L �b   �                            �L H                        8M �b                         lM H                        �M �b                         �M $H                        N �b                         :N 0H                        nN �b                         �N <H                        �N �b                         O HH                        JO �b                         �O TH                        �O �b                         P `H                        <P �b                         oP lH                        �P �b                         �P xH                        4Q �b                         iQ �H                        �Q �b                         �Q �H                        8R �b                         lR �H                        �R �b                         �R �H                        S  c        �                       =S �H                        tS c                         �S �H                        �S c                         T �H                        >T c                         nT �H                        �T  c                         �T �H                        @U $c                         �U �H                        �U 0c                         V �H                        FV @c     '                   �V I                        �V hc                         W I                        ZW tc                        �W  I                        �W �c                        5X ,I                        ~X �c                         �X 8I                        �X �c                         Y DI                        VY �c                         �Y PI                        �Y �d	                �                �Y ��                         �Y �d	         �Y �X	         Z �.          8Z �O	         nZ @K	         �Z �N                        �Z @O	         �Z �O	         �Z �e	         [ �e	         %[ pe	         8[ 0Y	         S[ `Z	     .text   �                       .data                           .bss    P                            n[ �d	    �                    �[ �c                          �[ \I                         �[ �X	                        �[ �c                          �[ hI                         \ �O	    ;                    S\ �c                          �\ tI                     .rdata       U                     �\ @K	    �                   �\ �c                          ] �I                         D] @O	    T                    w] d     -                    �] �I                         �] �O	    A                  �        ^ 4d                          :^ �I                         h^ �e	    W                    �^ @d                          �^ �I                         �^ pe	                        �^ Hd                          �^ �I                         _ 0Y	    0                   #_ Pd                          E_ �I                         g_ `Z	    �                   �_ `d                          �_ �I                         �_ �.                          �_ P$                          $` @$                          L` �\                          g` �\                          �` �\                          �`  ]                          �` �\                          �` P\                          �` @]                          a p\                          (a `\                          Ca �]                          ba p]                          �a P]�                                �a 0]                          �a  \                          �a �]                          b @\                          %b  ^                          Fb �]                          eb `]                          �b �]                          �b �]                          �b �]                          �b 0\                          c ]                          #c �\                          >c �\                          Zc �]                          zc �\                          �c  ]                          �c �\                          �c �]                          �c �    5                   �c �                          d p^     P                   d  ^     P                   -d 0    I                   =d 0         Gd  �    5                   |d  �         �d �a     P                   �d �a     �      P                   De ��    I                   ye ��         �e �	    4                   �e �	         f ��	    <                   0f ��	         Bf ��	    4                   Xf ��	         hf P�	    <                   �f P�	         �f P�	    Q                   �f P�	         g ��	    J                   g ��	         ,g ��	    Q                   ig ��	         �g ��	    J                   �g ��	         h �	                        8h �	         Zh �    �                   �h �         �h      �   	                �h           .i `�     x   	                <i �    K                    Li �         Vi �    �                   fi �         pi      �   	                �i           �i     �                   �i          �i �     $                  �i �          �i     �                   �i �               �i 0     �                   �i 0          j  �	                        0j  �	         Rj ��    �                   �j ��         �j ��    �   	                6k ��         ~k ��     x   	                �k `�    K                    �k `�         l 0�    �                   Jl 0�         yl ��    �   	                �l ��         �l ��    �                   m ��         Gm ��    ,                  m ��         �m ��    �                   �m ��         n ��    �                   Vn ��         �n ��                         �n �q     8                   �n `�     (                    �n pv     8                   o �     8                   o @�     8               .text   �                       .data                           .bss    P                            No ld                         _o �I     �                         po pd                         �o �I                        �o xd                         �o �I                        �o |d                         4p �I                        jp �d                         �p J                        �p �d                         �p J                        q �d                         +q J                        Bq �d                         �q (J                        �q �d                         �q 4J                        �q �d                         r @J                        r �d                         \r LJ                        �r �d                         �r XJ                        s �d                         ;s dJ                        ds �d     !                   �s pJ                        �s �d     (                   t |J         �                     Ht e                         Yt �J                        jt e     !                   {t �J                        �t ,e     $                   �t �J                        �t Pe                         �t �J                        �t `e     #                   �t �J                        �t �e                        u �J                         u �e                        6u �J                        Lu �e                         uu �J                        �u �e     !                   �u �J                        <v �e     )                   �v �J                        �v f                         w  K                        Fw f     !                   |w K                        �w 0f     $                   �w K                        x Tf                         Wx $K                 �             �x df     #                   �x 0K                        y �f                        ;y <K                        ty �f                        �y HK                        L�                               �y �:    )                   �y �:         z ��     P                   z �:    >                   $z �:         .z  �    )                   bz  �         �z �     P                   �z ��    >                   �z ��         ${ @�	    0                   <{ @�	         N{ ��	    0                   �{ ��	         �{ ��	    F                   �{ ��	         2| ��	    F                   J| ��	         \| P:    &                   �| P:         �| P8    �                   �| P8         0}  ;                        @}  ;         J}  <                        a}  <         r} 0<                        �      �} 0<         �} <                        �} <         ~ ��                        ,~ ��         <~ �0    �                   T~ �0         f~ �:    %                   v~ �:         �~  9    �                   �~  9         �~ �9    �                   �~ �9         �~ @7    
                  �~ @7         �~ @;    �                   �~ @;         �~ p    �                   	 p          �.    E                  2 �.         F P,    E                  ` P,         t `?    �                  � `?         � �=    S                  � �=         � P<    '                  � P<         � p                      (� p         4� 0    ;                  G� 0         T� �    B                  i� �         x� @    �                   �� @         �� �    �         �               Հ �         
�      w                   D�           x� P%    �                   �� P%         �� �    �                   �� �         �� �    �                   с �         ��  6                       ��  6         � �4    $                  "� �4         2� 0$                      F� 0$         T� 0     �                   g� 0          t� @#    �                   �� @#         �� !                      �� !         ʂ 0"                      � 0"         � ��                        %� ��         8�  �	    �                   w�  �	         �� ��	    �                   � ��	         .� P�	                       k� P�	         �� @�	                       ߄ @�	         � 0�	                       S� 0�	         ��  �	                       ǅ  �	         �� P�	    ~ �                        L� P�	         �� ��	                        � ��	         *� ��	                        z� ��	         ć �	    :                    � �	         P� ��	                        �� ��	         � ��	                        .� ��	         n� P    C                  �� P         �� �@                       �� �@         ȉ `    C                  � `         � 0?                       � 0?         "� �    C                  D� �         `� @?                       q� @?         |�      C                  ��           �� P?                       ˊ P?         ֊  	    C                  ��  	         � �=                       %� �=         0� �    C                  R� �         n�  A                       �  A         �� �    C                  �� �         ȋ A�                             ً A         �     C                  �          "� �=                       3� �=         >� p
    C                  `� p
         |� �=                       �� �=         �� �    C                  �� �         ֌ �=                       � �=         � �    C                  � �         2� �=                       D� �=         P� `�    &                   �� `�         � P�    �                   1� P�         x� 0�                        �� 0�         ڎ �                        � �         N� @�                        �� @�         ��  �                        %�  �         d� ;                        �� ;         Ґ �    N                   � �         D� ��    %                   x� ��         �� �    �                   ڑ �     �          � ��    �                   ?� ��         p� 0�                      �� 0�         ؒ P�    �                   � P�         @� @�    �                   z� @�         �� �    �                  � �         &� �    �                  e� �         �� p�    �                  Ӕ p�         � �    S                  7� �         f� `�    '                  �� `�         �� 0�    !                  0� 0�         `� ��    5                  �� ��         Ȗ �}    Y                  � �}         4� 0}    N                   l� 0}         �� 0�    �                  � 0�         8� �    F                   �� �         И 0�                       	� 0�         <� `�    �                   s� `�         �� P�    �                   ݙ P�         � �    1                  M� �      �         �� ��    "                  �� ��         �  �    #                  *�  �         \�  �    �                   ��  �         ě �    �                   �� �         .� ��                      o� ��         ��  �                      �  �         4�  ;                        q�  ;         �� �	    �                   � �	          � `�	                      b� `�	         �� ��	    �                  �� ��	         � 0�	    W                   j� 0�	         �� p�	                         � p�	         H� ��	                        �� ��	         � ��	    :                    +� ��	         n� ��	                        �� ��	         � ��	                        L� ��	         �� @y    D                  Ӣ @y         �  �                       I�  �         x� Pu    D            �            �� Pu          � @�                       5� @�         d� �v    D                  �� �v         � P�                       !� P�         P� �w    D                  �� �w         إ `�                       � `�         <� p    D                  �� p         Ħ ��                       �� ��         (� �z    D                  o� �z         �� �                       � �         � �{    D                  [� �{         ��  �                       Ѩ  �          �  t    D                  G�  t         �� У                       �� У         � `q    D                  3� `q         t� ��                       �� ��         ت �r    D                  � �r         `� ��                       �� ��         ī �n    D                  � �n         N� ��        �                     �� ��         �� Д                         ¬ �q     (                   Ь  �     '                    � �u     (                   4�  �                        B� �                    .text   �                       .data                           .bss    P                            t� �f                         �� TK                        �� �f                         �� `K                        �� �f                         � lK                        "� �f                         W� xK                        �� �f                         �� �K                        �� �f                         �� �K                        8� �f                         u� �K                        �� �f                         ˯ �K                        � �f                         � �K                        V� �f   �                           �� �K                        Ȱ g                         ٰ �K                        � g                         � �K                        � g                         R� �K                        �� g                         �� �K                        α $g                         � �K                        �� (g                         � L                        .� 4g                         ?� L                        P� 8g                        a�  L                        r� Xg                         �� ,L                        �� dg     #                   �� 8L                        �� �g                        Ѳ DL                        � �g                        �� PL                        � �g     L                   +� \L                        F� h     L   �                      a� hL                        |� Ph     T                   �� tL                        �� �h     T                   �� �L                        ĳ �h     D                   �� �L                        6� <i     D                   I� �L                        \� �i     H                   p� �L                        �� �i     L                   �� �L                        �� j                         Ŵ �L                        ڴ  j     L                   � �L                        R� lj                         �� �L                        ȵ xj     H                   ޵ �L                        �� �j     @                   � �L                        �  k     D                   2� �L                        H� Dk     P                   b� M                        |� �k     L          �               �� M                        �� �k     H                   �� M                        Զ (l     @                   � (M                        �� hl     D                   � 4M                        &� �l     H                   D� @M                        b� �l     H                   �� LM                        �� <m                         Ʒ XM                        � @m                         � dM                        `� `m     L                   �� pM                        � �m                         $� |M                        b� �m                         �� �M                        ޹ �m                         � �M                        Z� �m                         �� �M                        ֺ �m                         %� �M                        t� �m                       �        û �M                        � �m                         c� �M                        �� �m                         �� �M                        H� �m                         �� �M                        � �m                         /� �M                        v� �m     T                   �� �M                        �� 4n                         ξ  N                        � 8n     T                   � N                        &� �n                         8� N                        J� �n     T                   m� $N                        �� �n                         �� 0N                        �� �n     T                   ׿ <N                        �� <o                         � HN                        � @o     T                   A� TN                        d� �o                         v� `N�                              �� �o     T                   �� lN                        �� �o                         �� xN                        �� �o     T                   � �N                        8� Dp                         J� �N                        \� Hp     T                   � �N                        �� �p                         �� �N                        �� �p     T                   �� �N                        � �p                         � �N                        0� �p     T                   S� �N                        v� Lq                         �� �N                        �� Pq     T                   �� �N                        �� �q                         �� �N                        � �q                         V� �N                        �� �q                        �� O     �                         @� �q                         u� O                        �� �q                         ��  O                        &� �q                         s� ,O                        �� �q                         � 8O                        L� �q                         �� DO                        �� �q                         �� PO                        <� �q                         q� \O                        �� �q                        �� hO                        � r                         H� tO                        �� $r     #                   �� �O                        �� Hr                        (� �O                        `� `r                        �� �O                        �� xr     L                   � �O                        V� �r     L                   �� �O           �                   �� s     T                   � �O                        B� ds     T                   x� �O                        �� �s     D                   �� �O                        J� �s     @                   �� �O                        �� <t     H                   �� �O                        (� �t     L                   b� �O                        �� �t                         �� P                        � �t     X                   _� P                        �� 4u                          � P                        P� @u     H                   �� (P                        �� �u     <                   �� 4P                        4� �u     D                   n� @P                        �� v     L                   �� LP                        $� Tv     H                   _� XP                  �            �� �v     D                   �� dP                        � �v     @                   D� pP                        |�  w     D                   �� |P                        �� dw     H                   0� �P                        r� �w     H                   �� �P                        � �w                         B� �P                        �� �w                        �� �P                         � x     L                   C� �P                        �� dx     l                   �� �P                        � �x                         [� �P                        �� �x                         �� �P                        H� �x                         �� �P                        �� �x                         4� �P                        ~� �x                         ��  Q                        ��       �x                         e� Q                        �� �x     T                   �� Q                        <� Dy                         r� $Q                        �� Hy     T                   �� 0Q                        8� �y                         n� <Q                        �� �y     T                   �� HQ                        4� �y                         j� TQ                        �� �y     T                   �� `Q                        0� Lz                         f� lQ                        �� Pz     T                   �� xQ                        ,� �z                         b� �Q                        �� �z     T                   �� �Q                        (� �z                         ^� �Q                        ��  {     T                   �� �Q                        $� T{   �                            Z� �Q                        �� X{     T                   �� �Q                         � �{                         V� �Q                        �� �{     T                   �� �Q                        � |                         R� �Q                        �� |     T                   �� �Q                        � \|                         N� �Q                        �� `|     T                   �� R                        � �|                         M� R                        } p                         L�                               ��              �� �    	                    �� �         ��      	                    �           H� �                        z� �         �� �                         �� �          � �                         3� �          ^� �    	   �                       �� �         �� `    	                    �� `         "� �                        T� �         �� �                        �� �         �� �                        � �         8� 0P                       b� 0P         �� �     h                   ��  T                       ��  T         �� ��     h                   $� �    	                    Q� �         x� �    	                    �� �         �� p/                       �� p/         � ��     H                   0� �                        �� �         �� �                        � �         2� �                        V� �         t� `�    "                    �� `�         �Q               'Q               �� Ѕ	                       � Ѕ	         H� p�     0                   �� ��	                       �� ��	 �              � ��     0                   �f               b� 0I	                       �� 0I	         �� ��     x                   /� PJ	                       v� PJ	         �� ��     `                   �� H                       "� H         B� ��                         f�  r	                       ��  r	         �� p�     (                   6�  q	                       ~�  q	         �� ��     P   	                � �5                       V� �5         �� 4                       �� 4         iR               �Q               :�  P    $                   d�  P         �� �S    $                   �� �S         �� ��	    $                   � ��	         b� ��	    $                   �� ��	         Kg               �� @/    $                   � @/         0�  I	    $                   w�  I	         ��  J	    $ �                        ��  J	         @� �G    $                   f� �G         �� �q	    $                   �� �q	         � �p	    $                   X� �p	         �� �5    $                   �� �5         4� �3    $                   �� �3         >�              �� ��    #                   �� ��         &� p    #                   X� p         �� �    #                   �� �         �� �    #                   � �         H� 0    #                   w� 0         �� �    #                   �� �         �� 0    #                   2� 0         `�      #                   ��           �� �    #                   �� �         �     #                   4�          V� @    #                   � @         �� `g	    (                   �� `g	         �� ��     8                   �� 0g�      	    0                   
� 0g	          � �F	    (                   ;� �F	         P�  �     8                   i� �F	    0                   �� �F	         �� P)    (                   �� P)         ��  )    0                   ��  )         � �    (                   @� �         ]� P    0                   �� P         �� ��    T                   �� ��         �� p�                         �� `�                       � `�         /� �                       T� �         s� ��     X   
                �� p    $                   �� p         4� �B         �� �T         �� p�    �                  '� p�         N�  �    1  	                �  �         ��              ��              ��  a    s                   ��  a         �� �`    s                   %  �`         J  0b    ]               �          u  0b         �  �g    s                   �  �g         �  pg    s                    pg         :  i    ]                   e  i         � ��    L                   � ��         � ��     h                   � ��    L                    ��         +  �    H                   l  �         � �    H                   � �         # P�    G                   K P�         m `�    G                   � `�         � P     #                   � P           @    #                   D @         o 0    N                   � 0         � ��    N                   � ��          �     N                   H �          s �     N                   � �          �       #                   �            ' p�    #                   U p�         } @�    #                   � �      @�         � `�    L                   � `�           �     h                   4 p�    L                   W p�         t ��    H                   � ��         � Ј    H                   1 Ј         l �    G                   � �         �  �    G                   �  �          	 �    #                   1	 �         \	 �    #                   �	 �         �	 p    N                   �	 p         
 �    N                   7
 �         `
 0    N                   �
 0         �
 �    N                   �
 �          `    #                   G `         p �    #                   � �         � �    #                   � �          @N    �                   I @N         p �L    �                   � �L         �  O    �                   �  O    �            `M    �                   H `M         p @P                       � @P         � R    �                   � R          PP    �                   ? PP         f �R    �                   � �R         � 0Q    �                   � 0Q          T                       < T         ` ��	                       � ��	         � `�	                       5 `�	         x ��    k                    � ��         T 0�    k                    � 0�         2 ��	                       { ��	         � ��	                        ��	         J ��	                       � ��	         � �    ^                    3 �         � ��    S                    � ��         D  �	                       �  �	         � 0<    W                   � 0<          �;    W                   9�       �;         X  =    R                   }  =         � Pl	    I                   � Pl	         � 0�     H                   � `k	    I                    `k	          �k	    E                   N �k	         | �j	    E                   � �j	         �  l	    G                   �  l	          k	    G                   2 k	         J p    #                   t p         � �    #                   � �         � �    N                   
 �         ( @    N                   L @         j �    N                   � �         � �-    �                   � �-         � �+    �                    �+         > `.    �                   f `.         � �,    �                   � �,         � �/                       � �/          �H	                       [ �H	                � �H	                       � �H	         $ `)    _                    � `)         � �*    _                    h �*         � �)    _                    > �)         �  *    _                      *         |  )    _                    �  )         T  @I	                       �  @I	         �   J	                       #!  J	         d! �I	                       �! �I	         �!  �    ;                    F"  �         �" `�    >                    �" `�         H# ��    M                    �# ��         �# ��    <                    R$ ��         �$ `J	                       �$ `J	         0%  �    U                   P%  �         j% p�    U                   �% p�         �% И    Q                   �% И         & @�    Q                   I& @�         |& 0�    �                         �& 0�         �& ��    �                   �& ��         ' P                        7' P         d' p                        �' p         �' �                        �' �         .( @                        `( @         �( �                        �( �         �( P    B                    ) P         *) �    Q                    a) �         �) �    �                    �) �         �)     �                    *          P* ��    T                   p* ��         �* �E    �                  �* �E         �* �C    �                  �* �C         +  H                       <+  H         \+ �q	                       �+ �q	         �+ �q	                       ., �q	         p, �}    Z                    �, �}         ,- 0r	                       t- 0r	         �- `5                             	. `5         V. ��     (                   �.  5                       �.  5         D/ �5                       �/ �5         �/ @5                       :0 @5         �0  6                       �0  6         "1 �p	                       j1 �p	         �1 �p	                       �1 �p	         62 �    #                   �2 �         �2 @F    _                    L3 @F         �3 �E    _                    24 �E         �4 P    _                    5 P         �5 �    _                    6 �         �6 �F    _                    �6 �F         h7 q	                       �7 q	         �7 �3                       E8 �3         �8 0�     P   	                �8 `3                       39 `3         �9 �3                       �9 �3         ": �3                       v: �3               �:  4                       ;  4         ^; �f	    B                   z; �f	         �; @f	    B                   �; @f	         �; �f	    B                   �; �f	         �; �e	    B                   < �e	         :< �    #                   h< �         �<      #                   �<           �< �    ,                    = �         0= P                       Q= P         l= �g	    (                   �= �g	         �= �                        �= �         �= �    "                   .> �         Z> `(    �   
                �> `(         �> �     8                   �> �'    �   
                �> �'         ? )                       4? )         V? P(                       ~? P(         �? �)    (                   �? �)         �? ��         @ ��          @ �    �                         H@ �         j@ �    �                   �@ �         �@ �    �                   �@ �          A �    �                   )A �         LA �                       qA �         �A 0F	    B                   �A 0F	         �A �E	    B                   �A �E	         �A �E	    6                   B �E	         $B `E	    6                   AB `E	         XB P�                        �B P�         �B ��                        �B ��         �B  �    #                   C  �         :C �F	    (                   UC �F	         jC �    �                   �C �         �C `�     8                   �C �
    �                   �C �
         D p    �                   >D p         _D �    �                   �D �         �D �    (                   �D �         �D p�	    V                         E p�	         CE �z    �                  �E �z         F      9                  �F           �F �    �                  wG �         �G 0�	    V                    H 0�	         OH  ~                        jH ��	    V                   �H ��	         �H �#                         �H @~                        �H ��	    V                   2I ��	         `I �$                         |I �                        �I �7    �  #                �I �7         �I p�	    V                   [J p�	         �J  $                         �J �~                        @K ��	    V                   �K ��	         �K  $                         ?L �~                        �L ��	    V                   �L ��	         �L                           M �r     8                   8M �b    �  *                tM �b         �M       0�	    V                   �M 0�	         N                          =N �r     8                   ^N �[    �  *                �N �[         �N ��	    V                   1O ��	         �O  %                         �O `�                        P 0�	    V                   }P 0�	         �P �$                         !Q  �                        hQ ��	    V                   �Q ��	         �Q P                         �Q �s                        R  ~    d                  tR  ~         �R p�	    V                   2S p�	         �S �$                         �S p�                        T ��	    V                   zT ��	         �T �$                         U �     8                   bU 0�	    V                   �U 0�	         �U `$                         �U 0     8                   �U Я	    Q                         (V Я	         PV ��	    Q                   �V ��	         �V P�	    Q                   �V P�	         W P�	    Q                   9W P�	         dW в	    Q                   �W в	         X �	    Q                   rX �	         �X P�	    Q                    Y P�	         2Y P�	    Q                   �Y P�	         �Y ��	    Q                   FZ ��	         �Z �	    Q                   �Z �	         [ е	    Q                   _[ е	         �[ �	    Q                   \ �	         j\ ��	    Q                   �\ ��	         �\  �	    �                   �\  �	         &] @�    �                   �] @�         �] p�    L                   S^ p�         �^ ��    �  +                &_ ��         �_ �    �  +                �_ �         d` ��    M                  �` ��         a @�    ^                         �a @�         �a  {    �                  !b  {         ^b p�    <                   �b p�         c ��	    �                    Vc ��	         �c ��	    �                    �c ��	         �c �                      Ed �         �d `                      �d `         k              e ��    L                  ze ��         �e ��    6                   =f ��         �f ��    [                   �f ��         Bg @�    �                  �g @�         �g �    �                  bh �         �h  �    6                   %i  �         |i P�    [                   �i P�         *j  �    L                  �j  �         �j @�    8                   Yk @�         �k ��    [                   
l ��         ^l P�    �                  �l P�         0m ��    8                   �m ��  	             �m ��    �                   Cn ��         �n �    [                   �n �         Jo  �    S                  �o  �         "p �    H                   p �         �p `�    s                  Eq `�         �q `�    Q                   r `�         �              br �    �                  �r �         ^s �7    �                  �s �7         lt `                      �t `         `u �                      �u �         Xv �"    �  $                �v �"         `w P    7                  �w P         Nx     7                  �x          <y �C                      �y �C         "z �A                      �z �A         { �!    E  '                { �!         �{ �3    �                  g| �3         �| �5    �                  C} �5         �} �7    n  
      	                ~ �7         �~ `�    �                   `�         � p9    [                   � p9         b� `+    |                   Ѐ `+         8� �.                      �� �.         � �    s                  �� �         � 0:    [                   �� 0:         � `,    |                   Z� `,          ��    s                  C� ��         �� 9    [                   /� 9         �� �*    |                   � �*         p� P�    s                  � P�         l� �9    [                   ݈ �9         H� �+    |                   �� �+         � P    �	                  �� P         � �:    [                   �� �:         �� �,    |                   d� �,         ̌ �    �                  M� �         ȍ �:    [                   9� �:         �� �-          �                   � �-         �� `-    |                   �� `-         X� @�    �
  '                ڐ @�         V� `�    �
  (                ؑ `�         T�  �    [                  Ȓ  �         6� �                      �� �         � 0;    c                  �� 0;         � `�	         0� �                         U� �                         z�                          ŕ 0                         � �                         .� P                         w� p                         ��                          � �                         ,� �                         v� �                         �� 0                         �� ��                         ʗ `�                         � 0w                        � �                         &� ��                         H� �w                              j� ��     :                    ��  �     :                    �� ��                         � 0y                        <� ��                         Z� @�                         {�  �                         �� ��                         �� ��     !                    � �|     8                   � `�                         )�  �                         L� �v                        o�  �                         �� py                        ��  �                         � �y                        � ��     <                    V� @�     <                    �� ��     ;                    � ��     C                    1� px                        �  �     ;                    Ŝ ��     C                    � 0x                        a� @�                         �� �w                        ��  �                               ͝ �{     8                   �� ��     X                   !�  �     �                   I� �W                         v� �W                         �� `W                         ɞ PW                     .text   �                       .data                           .bss    P                            � �|                         $�  R                        Y� �|                         �� ,R                        ß �|                         �� 8R                        )� �|                         [� DR                        �� �|                         �� PR                        � �|                         &� \R                        [� �|                         �� hR                        š �|                         �� tR                        +� �|                         ]� �R                              �� �|                         �� �R                        � �|                         � �R                        I� �|                         t� �R                        �� �|                         ͣ �R                        �� �|                         )� �R                        W� �|                         |� �R                        �� �|                         �� �R                        O� �|                         �� �R                        �� �|                         إ �R                        ��  }                         %� �R                        M� }                         �� S                        � }                         +� S                        u� }                         �� S                        � }                         M� (S                        ��       }                         �� 4S                        � }                         ,� @S                        u� }                         �� LS                        �  }                         X� XS                        �� $}                         �� dS                        K� (}                         v� pS                        �� 0}                         ̫ |S                        �� 8}                         A� �S                        �� @}                         լ �S                        � H}                         D� �S                        i� P}                         �� �S                        �� X}                         A� �S                        �� `}                         �� �S                        ׮ h}                          � �S                        i� p}                               �� �S                        �� x}                         L� �S                        �� �}                         � �S                        ?� �}                         o�  T                        �� �}                         ұ T                        � �}                         :� T                        o� �}                         �� $T                        ٲ �}                         	� 0T                        9� �}                         l� <T                        �� �}                         Գ HT                        	� �}                         >� TT                        s� �}                         �� `T                        Ŵ �}                         � lT                        � �}                         A� xT                        k� �}                              �� �T                        �� �}                        µ �T                        ߵ  ~                        �� �T                        � ~                        3� �T                        O�  ~                        t� �T                        �� 0~                        �� �T                        � @~                        � �T                        +� P~                        O� �T                        s� `~                        �� �T                        �� t~                         ַ �T                        �� |~                         � �T                        C� �~                         i� U                        2A �B    G                     zA �~                          �A U                         �� �T    @                    �� �~                                ܸ  U                         � �~     T                   1� ,U                        _� �~     .                   �� 8U                    .rdata  p     �  M                 ù                           � DU                        � $                         G� PU                        s� (                         �� \U                        ˺ 0                         �� hU                        #� 4                         O� tU                        {� 8                         �� �U                        ӻ @                        �� �U                        � \                        ?� �U                        c� x                        �� �U                        � �                        )� �U                        k� �                        �� �U                              �� �                        � �U                        � �                         A� �U                        s� �                         �� �U                        ׾ �                         � �U                        /� �                         _� �U                        ��  �                         �� V                        � �                         %� V                        W� �                         �� V                        �� �                         �� (V                        � �                         D� 4V                        s� �                        �� @V                        �� 8�                        �� LV                        � T�                        E� XV                        �� p�                        �� dV                        � ��                              4� pV                        ]� ��                        �� |V                        �� Ā                         �� �V                        � Ȁ                         E� �V                        w� ̀                         �� �V                        �� Ԁ                         �� �V                        /� ܀                         a� �V                        �� �                         �� �V                        �� �                         '� �V                        W� ��                         �� �V                        �� �                         �� �V                        � ��     (                   A� �V                        o�  �     (                   ��  W                        �� H�     (                   �� W                        )� p�     (                         X� W                        �� ��                         �� $W                        �� ��     (                   � 0W                        9� ā     (                   g� <W                        �� �     (                   �� HW                        �� �     (                   "� TW                        Q� <�                         |� `W                        �� @�                         �� lW                        ;� D�                         �� xW                        �� H�                         A� �W                        �� P�                         &� �W                        �� X�                         �� �W                        -� \�                         w� �W                        �� `�                         � �W                        U� d�                               �� �W                        � l�                         r� �W                        �� t�                         � �W                        g� x�                         �� �W                        �� |�                         �� �W                        �� ��                         %� �W                        K� ��                        h� X                        �� ��                        �� X                        �� ��                        ��  X                        )� ܂                        ^� ,X                        �� ��                        �� 8X                        �� �                        �� DX                        � 0�                         :� PX                        e� 4�                         �� \X                        �� 8�                               �� hX                        � @�                         *� tX                        O� H�                         u� �X                        �� P�     (                   �� �X                        �� x�     (                   � �X                        ;� ��     (                   d� �X                        �� ȃ     (                   �� �X                        �� ��                         � �X                        )� �                         q� �X                        �� ��                         � �X                        I� ��                         �� �X                        '� �                         �� �X                        � �                         t� �X                        �� �                         R� Y                        �� �                         1�       Y                        �� $�                         �� Y                        1� (�                         y� (Y                        �� ,�                         	� 4Y                        Q� 0�                         �� @Y                        � 8�                         b� LY                        �� @�                         � XY                        s� H�                         �� dY                        -� P�                         u� pY                        �� T�                        �� |Y                        �� p�                         � �Y                        A� ��                        {� �Y                        �� ��                        �� �Y                        )� Ą     4                   O� �Y                        u� ��     4                   �� �Y                              �� ,�                         �� �Y                        )� 0�                         ]� �Y                        �� 4�                         �� �Y                        � 8�                         6� �Y                        i� <�                         �� �Y                        �� @�                         ��  Z                        � D�                         O� Z                        �� H�                         �� Z                        �� L�                         � $Z                        U� P�                        v� 0Z                        �� d�                         �� <Z                        �� h�                         � HZ                        3� l�                         Z� TZ                        �� p�                         �� `Z                              � t�                         \� lZ                        �� x�                         � xZ                        i� ��                         �� �Z                        �� ��                         O� �Z                        �� ��                         �� �Z                        K� ��                         �� �Z                        �� ��                         J� �Z                        �� ��                         �� �Z                        A� ��                         �� �Z                        �� ��                         � �Z                        e� ��                         �� �Z                        � ��                         �� �Z                        �� ��                         r� �Z                        �� ��                         d� [                              �� ��                         \� [                        �� ą                         P�  [                        �� ̅                         � ,[                        Y� Ѕ                         �� 8[                        � ԅ                         U� D[                        �� ؅                         �� P[                        S� ܅                         �� \[                        �� ��                         N� h[                        �� �                        �� t[                        ��  �                        �� �[                        � �                        5� �[                        W� 8�                        y� �[                        �� T�                         �� �[                        �� X�                         +� �[                              ]� \�                         �� �[                        �� d�                         �� �[                        �� h�                        
� �[                        '� x�                         Z� �[                        �� |�                         �� �[                        �� ��     &                   � �[                        C� ��     &                   k� \                        �� Ԇ                         �� \                        �� ؆                         � \                        7� ܆                        \� (\                        �� ��                        �� �                          �� 4\                         �� ��     &                   � @\                        D� �     &                   m� L\                        �� @�     &                   �� X\                              �� h�     &                   � d\                        >� ��                         d� p\                        �� ��                        �� |\                        �� ��                        �� �\                        �� ̇                           �\                        6  ԇ                         T  �\                        r  ܇                         �  �\                        �  ��                         �  �\                        " �                         G �\                        l �                        � �\                        � ��     (                   � �\                        � $�     (                    �\                        @ L�     (                   h �\                        � t�     (                   �  ]                              � ��                         ]                        ( ��                         Z ]                        � ��                         � $]                        X ̈                         � 0]                        V �                         � <]                        L ��                         � H]                        � �                         � T]                          �                         U `]                        � �     �                   � l]                        � ��                         X x]                        � ��                         	 �]                        x	 ��                         �	 �]                        �	 ��     �                   -
 �]                        j
 `�                         �
 �]                              �
 h�     �                    �]                        \ �                         � �]                          �                         � �]                        � $�                          �]                        V ,�                         � �]                          D�                         � �]                        � L�                         C �]                        � T�                         � ^                         \�                         = ^                        l d�                         �  ^                        � l�                          ,^                        4 t�                         f 8^                        � |�                         � D^                        R ��                         � P^                                ��                         E \^                        ~ ��                         � h^                        < ��                         � t^                        � ��                         0 �^                        f ��                         � �^                        " ��                         � �^                        � ��                          �^                        B ċ                         v �^                        � Ћ                          �^                        t ��                         � �^                        L �     |                   � �^                        * h�     |                   � �^                         �     :                   i �^                        �  �                         . �^                        � !      (�                         � _                         @�                         | _                        � L�                          _                        X T�                         � (_                        � \�     <                    4_                        b ��     <                   � @_                        � ԍ                         _  L_                        �  �                         *! X_                        �! �                         �! d_                        >" ��                         �" p_                        �" �                         g# |_                        �# 0�                         2$ �_                        �$ 8�                         �$ �_                        F% @�                         �% �_                         & X�     "                          ~& �_                        �& `�                         7' �_                        �' h�                         �' �_                        l( ��                         �( �_                        () ��                         �) �_                        �) ��                         C* �_                        �* ��                          + �_                        ~+ ��                         �+  `                        :, Ȏ                         �, `                        - �                         x- `                        �- �                         X. $`                        �. �                         e/ 0`                        �/ �                         n0 <`                        �0 4�                         l1 H`                        �1 L�          #                     t2 T`                        �2 d�                         w3 ``                        �3 |�                         m4 l`                        �4 ��                         _5 x`                        �5 ��                         J6 �`                        �6 ď     <                   <7 �`                        �7  �     /                   ,8 �`                        �8 0�     /                   9 �`                        �9 `�     +                   �9 �`                        f: ��     T                   �: �`                        j; ��                         �; �`                        N< �                         �< �`                        ,= �                         �= �`                        > �     J                   �> �`                        ? T�                  $             �? �`                        �? \�                         g@ a                        �@ d�     J                   XA a                        �A ��                         LB  a                        �B ��                         -C ,a                        �C ��     J                   D 8a                        �D �                         E Da                        �E �                         �E Pa                        bF �     T                   �F \a                        fG p�                         �G ha                        JH x�                         �H ta                        (I ��     S                   �I �a                        ,J Ԓ                         �J �a                        K ܒ                         �K �a                        �K �                         %      eL �a                        �L ��     6                   WM �a                        �M ,�     6                   ]N �a                        �N d�     4                   UO �a                        �O ��     4                   @P �a                        �P ̓                         .Q �a                        �Q `�	    �                    �Q �                          R �a                     .ctors  H�	                        L�                               \R �^    !                   lR �^         vR 0�     P                   �R `^    6                   �R `^         �R p�    !                   �R p�          S `�     P                   2S 0�    6                   fS 0�         �S ��	    (                   �S ��	         �S `�	    (                   �S `�	         0T p�	    >                   HT p�	 &              ZT  �	    >                   �T  �	         �T  ^                       U  ^         6U �[    �                   nU �[         �U �^                        �U �^         �U �_                        �U �_         �U �_                        V �_         JV �_                        kV �_         �V pI    K                   �V pI         �V C    �                   �V C         �V �E    �   
                �V �E         �V �C    �                   W �C         ,W �D    �                   PW �D         nW @^                       ~W @^         �W �\    �                   �W �\         �W  ^                        �W  ^         �W p\    i                   �W p\         �W �]    �                   �W �]         �W �Z    �                   X �Z         X �^    �                 '        ,X �^         8X pB    �                   MX pB         \X @H    o                   uX @H         �X �G    o                   �X �G         �X I    `                   �X I         �X �H    `                   �X �H         Y  `    V                  <Y  `         nY  A    A                  �Y  A         �Y �F    A                  �Y �F         �Y ��                        �Y ��         �Y �	    p                   !Z �	         \Z ��	                       �Z ��	         �Z Ш	                       [ Ш	         V[ ��	    ~                   �[ ��	         �[  �	                        :\  �	         �\ @�	                        �\ @�	         ] ��	    :                    e] ��	         �]  �	                        �]  �	         @^ `�	                        �^ `�	         �^ ��	    �       (                 _ ��	         h_ ��	                       �_ ��	         �_ ��	                       ` ��	         L` ��	                       �` ��	         �`  �	    P                   �`  �	         4a ��	    P                   ra ��	         �a P�	    P                   �a P�	          b @R                      ?b @R         Xb �a                       hb �a         rb �a    (                   �b �a         �b �a                       �b �a         �b `T                      �b `T         �b �a                       �b �a         �b  b                       c  b         c �a                       "c �a         ,c �K                      Kc �K         dc `a                       tc `a         ~c �V                      �c �V         �c 0b                       �c 0b         �c �X    )                        �c �X         d @b                       d @b         "d �M                      Ad �M         Zd pa                       jd pa         td �a    	                   �d �a         �d P    .                  �d P         �d �a                       �d �a         �d �I                      e �I         e �_                       .e �_         :e ��                       �e ��         �e p�    �                   f p�         bf ��                        �f ��         �f p�                        g p�         8g ��                        �g ��         �g ��                        h ��         Nh ��    K                   �h ��         �h 0�    �                   �h 0�         .i ��    �   
                fi ��         �i �    �                   �i �         j *      �    �                   \j �         �j �                       �j �          k ��    �                   4k ��         bk ��                        �k ��         �k  �    p                   @l  �         �l @�    �                   �l @�         �l p�    �                   %m p�         Vm ��    �                   �m ��         �m ��    �                   �m ��         ,n `�    o                   jn `�         �n �    o                   �n �         o 0�    `                   So 0�         �o Ю    `                   �o Ю         �o ��    V                  Ep ��         �p 0�    Q                  �p 0�         �p ��    A                  -q ��         bq 0;                        �q 0;         �q `�	    E                   r `�	         Rr ��	                       �r ��	    +           �r �	                       s �	         Ls  �	    W                   �s  �	         �s @�	                        0t @�	         xt ��	                        �t ��	         u ��	    :                    [u ��	         �u `�	                        �u `�	         6v ��	                        |v ��	         �v ��	    �                  w ��	         ^w  �	                       �w  �	         �w @�	    P                   x @�	         Zx `�	    I                   �x `�	         �x ��	    �                  y ��	         Ny 0�    �                  �y 0�         �y ��                       z ��         2z ��    (                   fz ��         �z ��                       �z ��         �z  �    �                  :{  �         x{ ��                       �{ ��         �{ ��                       |,       ��         <| ��                       p| ��         �| ��    �                  �| ��          } 0�                       T} 0�         �} к    �                  �} к         ~  �                       8~  �         f~ ��    �                  �~ ��         �~ �                        �         J ��    �                  � ��         � @�                        � @�         .� p�    	                   b� p�         �� P�    �                  Ԁ P�         � P�                       F� P�         t� �    �                  �� �         �� ��                       0� ��         `� ��                         n�  r     (                   |� `�     '                    �� �u     (                   �� 0�                        � �                    .text   �                   -          .data                           .bss    P                             � �                         1� �a                        B� �                         S� b                        d� ��                         �� b                        ΃ ��                         � b                        8�  �                         Q� (b                        j� �                         �� 4b                        � �                         �� @b                        � �                         S� Lb                        �� �                         Ʌ Xb                        � �                        ;� db                        t� <�                         �� pb                        �� @�                         �� |b                        Ɔ D�                         �� �b                        .      6� L�                         X� �b                        z� T�                         �� �b                        �� `�     <                   Ň �b                        ڇ ��     @                   � �b                        � ܔ     <                   "� �b                        @� �     <                   e� �b                        �� T�                         �� �b                        �� X�                        �� �b                        Έ x�                         � �b                        � |�                         �  c                        � ��                         -� c                        @� ��                        S� c                        f� ��                        y� $c                        �� ĕ                        �� 0c                        �� ؕ  /                             ҉ <c                        � ��                         � Hc                         � �                        8� Tc                        P� ��                        h� `c                        �� �     P                   �� lc                        � `�     P                   � xc                        � ��     T                   0� �c                        H� �                         b� �c                        |� �                         �� �c                         � �                         B� �c                        �� �                         ǌ �c                        
� �                         Y� �c                        �� ,�                         �� �c                        F� 0�                         �� �c                        � 4�      0                         2� �c                        |� 8�                         ̏ �c                        � <�                         c� �c                        �� @�     d                   �� d                        T� ��                         �� d                        Α ��                         �  d                        H� ��                         �� ,d                         ��                         � 8d                        @� ȗ                         � Dd                        �� ԗ                         �� Pd                        <� ��     d                   \� \d                        |� D�                         �� hd                        �� H�                         �� td                        �� L�                         є �d                        � P�     d        1                 � �d                        "� ��                         3� �d                        D� ��                         U� �d                        f� ��                         w� �d                        �� ��     d                   �� �d                        ȕ $�                         ٕ �d                        � (�     d                   
� �d                        *� ��                         ;� �d                        L� ��     d                   l� �d                        �� ��                         �� �d                        �� ��     d                   Ζ e                        � \�                         �� e                        � `�                         !� e                        2� d�     `                   R� (e                        r� Ě                     2          �� 4e                        �� ̚     d                   �� @e                        ؗ 0�                         � Le                        �� 4�                         L� Xe                        �� 8�                        � de                        6� X�                         k� pe                        �� \�                         ޙ |e                        � `�                         i� �e                        �� h�                         �� �e                        B� p�                         �� �e                        �� |�     <                   �� �e                        2� ��     @                   k� �e                        �� ��     <                   � �e                        (� 4�     <                   q� �e                        �� p�                         � 3      �e                        $� t�                        Y� �e                        �� ��                         ۞ �e                        (� ��                         u�  f                         ��                         �� f                        2� ��                        j� f                        �� ̜                        ڠ $f                        � ��                        M� 0f                        �� ��                         ǡ <f                        � ��                         E� Hf                        �� �                        �� Tf                        �� �                        8� `f                        t� ,�     P                   £ lf                        � |�     T                   G� xf                        ~� Н     T                   �� �f     4                         �� $�                         4� �f                        r� (�                         �� �f                        �� 0�                         8� �f                        z� 4�                         �� �f                         � 8�                         O� �f                        �� D�                         � �f                        <� H�                         �� �f                        ި L�                         (� �f                        r� P�                         © �f                        � T�                         Y� �f                        �� X�     d                   �� g                        J� ��                         �� g                        Ϋ Ğ                         �  g                        V� О                         �� ,g         5                     ֬ ؞     d                   � 8g                        Z� <�     `                   �� Dg                        � ��                         � Pg                        N� ��                         �� \g                        �� ��                         � hg                        "� ��     `                   g� tg                        �� �                         � �g                        � �                         K� �g                        �� �                         �� �g                        � �     `                   /� �g                        t� t�                         �� �g                        ޱ x�     `                   #� �g                        h� ؠ                         �� �g                        Ҳ ܠ     `                   � �g                 6             \� <�                         �� �g                        Ƴ @�     d                   � �g                        P� ��                         �� �g                        �� ��                         � h                        $� ��     `                   i� h                        �� �                         � h                        � �     `                   _� (h                        �� t�                         ݶ 4h                        } �                         � ��                          E� P�         i� ��     .text   �                       .data                           .bss    P                            �� ��    o                   ɷ x�                          � @h                     .rdata                             9� P�    �                    c� ��                          7      �� Lh                         �� ��                        � ��                          � Xh                         H� p                        �� p                          ʹ �                        � �         >� �                        �� �         �                          H�           �� P                        ѻ P         � P                        B� P         z� �                        �� �         �                         .�          f� �                        �� �         ڽ p                        � p         \� �                         �� �          о �#                        -� �#         �� �#                        ڿ �#         *� P                        c� P         �� @%                        �� @%         � �%                        J� �% 8              ��  %                        ��  %         �� �$                        5� �$         l�                         ��           �� �     �                   � '                       <� '         l� ��     �                   �� �    (                   �� �         � �&    (                   <� �&         l�     �                   ��          ��  #    �                    �  #         X�       M                   ��            �� 0    L                    � 0         4� 0    �                   q� 0         ��  "    �                   ��  "         � @                       R� @         �� �    n                   �� �         
� 0<                       F� 0<         |�      #                   ��           �� �    M                   W� �         ��      Q 9                        �           `� �    #                   �� �         �� `    #                   � `         F�      �                   ��           �� �    p                   �� �         &� �    +                   `� �         �� �                        �� �         � `    >                   D� `         |�      =                   ��           �� �    E                   (� �         \�                          ��           �� �    C                   � �         6�      C                   l�           �� �;                        �� �;         � �;                        F� �;         z�  <                        ��  <         �� `                        $� `         X� �                        �� �         ��  <                        �  <         B� �;:                              |� �;         �� <                        �� <          � �                        Z� �         �� �                        �� �         � �    k                   =� �         r� `                        �� `         �� p                        2� p         n� P    G                   �� P         �� �    G                   � �         J� `    N                   �� `         �� �    �                   �� �         *� ��	                       |� ��	         �� 0'                       �� 0'         .� �$    n                   u� �$         �� �<                       �� �<         (� %    #                   h� %         �� �    M                   � �         ^�      Q                   ��           � �#    #                   H� �#     ;          ~� P$    ,                   �� P$         ��  !    �                   -�  !         b� p     q                   �� p          �� �    +                   � �         @� �                        |� �         �� P%    >                   �� P%         (� $    @                   d� $         �� �    >                   �� �         �                          E�           |� �&    C                   �� �&         �� �%    C                   � �%         H� p<                        �� p<         �� P<                        �� P<         &� �<                        a� �<         �� `                        �� `         � �                        D� �         ~� �<                        �� �<         �� `<                        (� `<         \� �<                        �� <      �<         �� �                        � �         :� �                        w� �         �� �!    k                   �� �!         � `                        `� `         �� p                        �� p         � @&    G                   T� @&         �� �%    G                   �� �%         �� P'    N                   0� P'         d� �    �                   �� �         �� ��	                       (� ��	         t� ��     )                    �� �w                        ��  �     )                    � �w                    .text   �                       .data                           .bss    P                            D� ��                         �� dh                        �� ��                         � ph                        J� ��                         �� |h                  =            � Ģ                         ]� �h                        �� Ȣ                         �� �h                        (� ̢                         g� �h                        �� Т                         �� �h                        $� Ԣ                         c� �h                        �� آ                         �� �h                        � ܢ                         c� �h                        �� �                         �� �h                        $� �                         �� �h                        �� �                         7� �h                        �� �                         ��  i                        � �                         A� i                        �� ��                         �� i                        �� ��                         =� $i                        |�>       ��                         �� 0i                        ��  �                         /� <i                        f� �                         �� Hi                        �� �                         � Ti                        B� �                         y� `i                        �� �                         �� li                        .� ,�                         m� xi                        �� @�                         �� �i                        "� H�                         ]� �i                        �� P�                         �� �i                        � d�                         R� �i                        �� x�                         �� �i                        �� |�                         F� �i                        �� ��                         �� �i                        � ��   ?                            I� �i                        �� ��                         �� �i                        N� ��                         �� �i                        � ��                         A� �i                        ~� ��                         �� j                        �� ��                         6� j                        r� ȣ                         ��  j                        �� У                         %� ,j                        `� ԣ                         �� 8j                        �� أ                         � Dj                        X� ܣ                         �� Pj                        �� �                         � \j                        H� �                         �� hj                        �� �                         �� tj                        2 	 �        @                       i 	 �j                        � 	 �                         � 	 �j                        	 ��                         S	 �j                        �	 ��                         �	 �j                        	 ��                         A	 �j                        |	  �                         �	 �j                        �	 �                         :	 �j                        v	 �                         �	 �j                        �	 �                         (	 �j                        d	 �                         �	 �j                        �	 �                         	 �j                        V	 �                         �	 k                        �	  �                         	 k                        T	 $�                         �	 k                        �	 (�                A               	 (k                        P	 ,�                         �	 4k                        �	 0�                         	 @k                        <	 8�                         y	 Lk                        �	 D�                         			 Xk                        \		 L�                         �		 dk                        �		 P�                         
	 pk                        Z
	 p�                         �
	 |k                        �
	 x�                         	 �k                        V	 |�                         �	 �k                        	 ��                         u	 �k                        �	 ��                         	 �k                        J	 ��                         �	 �k                        �	 ��                         	 �k                        >	 ��                       B        z	 �k                        �	 ��                         �	 �k                        ,	 ��                         i	 �k                        �	 ��                         �	 �k                        $	 ��                         a	  l                        �	 ��                         �	 l                        	 ��                         R	 l                        �	 ��                         �	 $l                        �	 ��                         5	 0l                        l	 Ĥ                         �	 <l                        �	 Ȥ                         	 Hl                        Z	 ̤                         �	 Tl                        �	 Ф                         	 `l                        H	 Ԥ                         �	 ll                        �	 ؤ                         	 xlC                              B	 ܤ                         }	 �l                        �	 �                         �	 �l                        0	 �                         k	 �l                        �	 �                         �	 �l                        "	 �                         ^	 �l                        �	 ��                         �	 �l                         	 ��                         c	 �l                        �	 ��                         �	 �l                        	  �                         W	 �l                        �	 �                         �	 �l                        	 �                         E	 �l                        �	 �                         �	 m                        (	 ��                        o	 ��                          �	 `�                        �	 `�     D          :	 P�                        �	 P�         �	  �                        	  �         V	  �                        �	  �         �	 ��                        7	 ��         |	 0�                        �	 0�         	  �                        \	  �         �	 ��    m                   �	 ��         0 	 ��                       z 	 ��         � 	 ��                       !	 ��         L!	 н    �                   �!	 н         �!	 @�    	                   3"	 @�         �"	 0�                        �"	 0�         #	  �                        k#	  �         �#	 ��    (                   $	 ��         F$	 ��    (                   �$	 ��         �$	 А                        1%	 А         t%	 ��                        �%	 ��         
&	  �                       U&	  �         �&	  �                       �&	 E       �         *'	 ��    $                   u'	 ��         �'	 `�                       2(	 `�         �(	 @�                       )	 @�         �)	 ��                       �)	 ��         0*	 ��                       �*	 ��         �*	 `�                        +	 `�         b+	 @�    �                   �+	 @�         �+	 p�    ;                  A,	 p�         �,	 0�    `                   �,	 0�         -	 ��                        R-	 ��         �-	 ��                        �-	 ��         .	 @�                        J.	 @�         �.	 `�                        �.	 `�         
/	 ��                       P/	 ��         �/	 ��                       �/	 ��         0	 0�    K                    Y0	 0�         �0	 P�    K                    �0	 P�         1	 ��    `                    ^1	 ��         �1	 ��    `              F            �1	 ��         *2	 0�                       j2	 0�         �2	 �                       �2	 �         3	 0�                       b3	 0�         �3	 P�    �                   �3	 P�          4	 ��                        d4	 ��         �4	 p�                        �4	 p�         &5	 ��                        h5	 ��         �5	 @�                        �5	 @�         $6	 ��                        i6	 ��         �6	 ��                        �6	 ��         .7	 ��    
                    q7	 ��         �7	 P�    
                    �7	 P�         08	 ��                        v8	 ��         �8	 `�                        �8	 `�         89	 ��                        9	 ��         �9	 ��    
                    :	 ��         D:	 `�                        �:	 `�         �:	 ��                        ;	 ��         L;	  �         G                     �;	  �         �;	 ��                        <	 ��         `<	  �                      �<	  �         �<	 ��    I                   3=	 ��         z=	 ��                        �=	 ��         �=	 ��    	                    A>	 ��         �>	 �                        �>	 �         �>	 ��                        <?	 ��         v?	 �    %                   �?	 �         �?	 P�    %                   5@	 P�         p@	 P�                        �@	 P�         �@	 ��                        7A	 ��         vA	 ��                        �A	 ��         �A	 P�                        :B	 P�         xB	 `�    w                   �B	 `�         �B	 ��    i                   :C	 ��         |C	 ��                       �C	 ��         D	 ��    �                   PD	 ��         �D	 ��    _                   �D	 ��         E	 ��  H        *                   �E	 ��         �E	  �    T                   QF	  �         �F	 ��                       �F	 ��         @G	 �                      �G	 �         �G	 ��    !                   "H	 ��         bH	 ��    @                   �H	 ��         �H	 ��                       -I	 ��         lI	 @�                        �I	 @�         �I	 ��    )                   2J	 ��         lJ	  �    @                   �J	  �         �J	 `�    6                   `K	 `�         �K	 ��    H                   L	 ��         RL	 P�                       �L	 P�         .M	 ��    3                   �M	 ��         N	 ��    �                  QN	 ��         �N	 ��    M                   �N	 ��         *O	 ��                       rO	 ��         �O	 P�    (                   
P	 P�         ZP	  �                        �P	  �         I      
Q	 P�    1                   QQ	 P�         �Q	 ��    =                   �Q	 ��         "R	 ��    1                   dR	 ��         �R	 @�    @                   �R	 @�         .S	  �    <                   wS	  �         �S	 ��    J                   T	 ��         LT	  �    V                   �T	  �         .U	 @�    I                   �U	 @�         V	 ��    V                   �V	 ��         �V	 ��    V                   eW	 ��         �W	 ��    Y                   ZX	 ��         �X	 ��    u                   &Y	 ��         lY	 @�    �                   �Y	 @�         Z	 @�    V                   �Z	 @�         �Z	 ��    V                   m[	 ��         �[	 ��    D                   ]\	 ��         �\	 @�    h                   "]	 @�         f]	 ��    V                   �]	 ��         �]	 `�    q                   b^	 `� J              �^	 ��    �                   _	 ��         ^_	 ��                       �_	 ��         �_	 �                       .`	 �         l`	 ��    C                   �`	 ��         �`	 ��    -                   Da	 ��         �a	 `�    H                   �a	 `�         b	 ��    H                   Pb	 ��         �b	 @�    7                   �b	 @�         <c	  �    7                   �c	  �         �c	 p�    h                   )d	 p�         jd	 ��    �                    �d	 ��         �d	 ��                        5e	 ��         te	 ��                        �e	 ��         �e	 ��                        Df	 ��         �f	  �    �                   �f	  �         g	 ��                       _g	 ��         �g	 ��    0                   �g	 ��         *h	  �    B                   oh	  �         �h	 ��    m                 K        �h	 ��         :i	 `�                       �i	 `�         �i	 ��    0                   j	 ��         Rj	 p�    0                    �j	 p�         �j	 @�    r                   *k	 @�         vk	 ��                       �k	 ��         l	 �    0                   gl	 �         �l	 І                       m	 І         Jm	 @�    s                   �m	 @�         �m	 ��                       8n	 ��         �n	 �    0                   �n	 �         o	 Ѕ    0                    lo	 Ѕ         �o	 0�    r                   
p	 0�         Zp	 ��                       �p	 ��         q	  �    0                   Wq	  �         �q	 ��    D                    �q	 ��         Fr	 `�    [                   �r	 `�         �r	 ��                       @s	 ��         �s	 0�    0                   �s	 0�         2t	 Ї    0         L                 �t	 Ї         �t	 Ѝ    Q                   u	 Ѝ         `u	 P�    }                   �u	 P�         �u	 Џ    �                   Cv	 Џ         �v	 `�    b                   �v	 `�         w	 0�    �                   cw	 0�         �w	 Ў    ~                   �w	 Ў         :x	 ��                        �x	 ��         �x	 ��                        0y	 ��         ~y	 ��                        �y	 ��         z	 ��                        qz	 ��         �z	 ��	    �                   {	 ��	         b{	 ��	    �                   �{	 ��	         |	  �    �                   �|	  �         }	 ��                       �}	 ��         �}	  �                       n~	  �         �~	 `�    �                   l	 `�         �	 ��                       A�	 ��         ��	 ��                       ̀	 ��         �	 `�    M      �                   }�	 `�         �	 `�                       (�	 `�         f�	 ��                       ��	 ��         �	 `�	    \                   ;�	 `�	         ��	  �                       փ	  �         �	  �                       l�	  �         ��	 ��    �                   "�	 ��         ��	 ��    B                   ԅ	 ��         �	 ��    B                   b�	 ��         ��	 ��    L                   �	 ��         ,�	 �    L                   r�	 �         ��	 @�    L                   ��	 @�         B�	 `�    L                   ��	 `�         ҈	  �                       �	  �         \�	 @�                       ��	 @�         �	 ��    ?                   -�	 ��         n�	  �    ?                   ��	  �         ��	 ��                       Q�	 ��         ��	 ��                       �	 ��         V�	 N      ��                       ��	 ��         �	 �                       =�	 �         ��	 Ќ    w                   ͍	 Ќ         �	 ��    
                    ��	 ��         �	 ��    
                    b�	 ��         Џ	 �[                     .text   �                       .data                           .bss    P                            �	  �                         [�	 m                        ��	 $�                         �	  m                        5�	 (�                         }�	 ,m                        ő	 ,�                         �	 8m                        a�	 0�                         ��	 Dm                        ��	 4�                         K�	 Pm                        ��	 8�                         �	 \m                        3�	 <�                         ��	 hm                    .rdata  0     �              O            ͔	 @�                         �	 tm                        c�	 H�                         ��	 �m                        ��	 L�                         D�	 �m                        ��	 P�                         ݖ	 �m                        +�	 \�                         �	 �m                        ӗ	 `�                         $�	 �m                        u�	 d�                         ǘ	 �m                        �	 h�                         e�	 �m                        ��	 p�                         �	 �m                        [�	 x�                         ��	 �m                        �	 |�                         >�	 �m                        ��	 ��                         ٛ	 �m                        %�	 ��                         q�	 n                        ��	 ��                         	�	 n                        U�P      	 ��                         Ν	 n                        G�	 ��                         ��	 (n                        9�	 ��                         ��	 4n                        �	 ��                         8�	 @n                        ��	 ��                         ٠	 Ln                        %�	 ��                         r�	 Xn                        ��	 ��                         �	 dn                        [�	 ȥ                         ��	 pn                        �	 ԥ                         .�	 |n                        o�	 إ                         ��	 �n                        �	 ܥ                         6�	 �n                        {�	 �                         ��	 �n                        �	 �                         L�	 �n                        ��	 �                         ڥ	 �n                        !�	 �   Q                            e�	 �n                        ��	 �                         �	 �n                        1�	 ��                         z�	 �n                        ç	 ��                         �	 �n                        U�	 ��                         ��	 �n                        ר	  �                         �	  o                        Y�	 �                         ��	 o                        �	 �                        '�	 o                        k�	 �                         ��	 $o                        ��	  �                         ;�	 0o                        ��	 $�                         ī	 <o                        �	 (�                         K�	 Ho                        ��	 ,�                         լ	 To                        �	 0�                         b�	 `o                        ��	 4�        R                       �	 lo                        1�	 8�                         v�	 xo                        ��	 <�                         �	 �o                        I�	 @�                         ��	 �o                        ӯ	 D�                         �	 �o                        c�	 H�                         ��	 �o                        �	 L�                         4�	 �o                        y�	 P�                         ��	 �o                        �	 T�                         P�	 �o                        ��	 X�                         �	 �o                        +�	 \�                         r�	 �o                        ��	 l�                        �	 �o                        U�	 ��                         ��	 �o                        ߴ	 ��                         %�	 p                        k�	 ��                S               ��	 p                        �	 ��                         0�	  p                        q�	 ��                         ��	 ,p                        ��	 ��                         9�	 8p                        {�	 ��                         ��	 Dp                        �	 ��                         K�	 Pp                        ��	 ��                         ո	 \p                        �	 ��                         ^�	 hp                        ��	 ��                         �	 tp                        %�	 Ȧ                         n�	 �p                        ��	 ئ                         �	 �p                        K�	 �                        ��	 �p                        ݻ	 �                         #�	 �p                        i�	 ��                         Լ	 �p                        ?�	 �                       T        ��	 �p                        �	 �                         c�	 �p                        ��	 �                         ��	 �p                        O�	 $�                         ��	 �p                        ݿ	 ,�                         $�	 �p                        k�	 4�                         ��	 �p                        ��	 8�                         >�	 q                        ��	 @�                         ��	 q                        �	 H�                         O�	 q                        ��	 P�                         �	 (q                        q�	 \�                         ��	 4q                        �	 d�                         w�	 @q                        ��	 h�                         W�	 Lq                        ��	 t�                         �	 Xq                        e�	 ��                         ��	 dqU                              ��	 ��                         F�	 pq                        ��	 ��                         ��	 |q                        =�	 ��                         ��	 �q                        ��	 ��                         =�	 �q                        ��	 ��                         ��	 �q                        �	 ��                         `�	 �q                        ��	 ̧                         ��	 �q                        9�	 ԧ                         ��	 �q                        ��	 ܧ                         �	 �q                        g�	 �                         ��	 �q                        Q�	 �                         ��	 �q                        9�	 ��                         ��	 �q                        #�	 ��                         ��	  r                        �	 �                         ��	 r     V                         �	 �                         j�	 r                        ��	 �                         �	 $r                        U�	  �                         ��	 0r                        S�	 (�                         ��	 <r                        ?�	 0�                         ��	 Hr                        C�	 8�                         ��	 Tr                        ��	 H�                         "�	 `r                        k�	 T�                         ��	 lr                        Q�	 d�                         ��	 xr                        ��	 p�                         3�	 �r                        }�	 t�                         ��	 �r                        �	 x�                         S�	 �r                        ��	 ��                         ��	 �r                        1�	 ��                         y�	 �r           W                   ��	 ��                         �	 �r                        G�	 ��                         ��	 �r                        ��	 ��                         V�	 �r                        ��	 ��                         ��	 �r                        =�	 ��                         ��	 �r                        ��	 ��                         �	 �r                        W�	 ��                         ��	 s                        ��	 Ĩ                         0�	 s                        �	 Ȩ                         ��	  s                        �	 ܨ                         [�	 ,s                        ��	 �                         ��	 8s                        5�	 �                         {�	 Ds                        ��	 ��                         �	 Ps                        U�	 �                         ��	 \s                  X            ��	 �                         4�	 hs                        }�	 �                         ��	 ts                        �	 �                         ^�	 �s                        ��	 ,�                         �	 �s                        Y�	 0�                         ��	 �s                        ��	 <�                         M�	 �s                        ��	 @�                         ��	 �s                        A�	 P�                         ��	 �s                        ��	 T�                         8�	 �s                        ��	 `�                         ��	 �s                        '�	 d�                         ~�	 �s                        ��	 t�                         -�	 �s                        ��	 x�                         ��	 �s                        1�	 ��                         ��	 t                        ��Y      	 ��                         /�	 t                        ��	 ��                         ��	 t                        3�	 ��                         ��	 (t                        ��	 ��                         0�	 4t                        ��	 ��                         ��	 @t                        �	 ��                         i�	 Lt                        ��	 ĩ                         �	 Xt                        W�	 Щ                         ��	 dt                        ��	 �                         7�	 pt                        ��	 �                         ��	 |t                        �	 ��                         r�	 �t                        ��	  �                         �	 �t                        q�	 �                         ��	 �t                        �	 �                         m�	 �t                        ��	 �   Z        "                   �	 �t                        m�	 0�                         ��	 �t                        �	 P�                         ��	 �t                        9�	 \�                         ��	 �t                        �	 `�                         ��	 �t                        �	 d�                         ��	 �t                        +�	 p�                         u�	  u                        ��	 t�                         	�	 u                        S�	 x�                         ��	 u                        /�	 ��                         t�	 $u                        ��	 ��                         ��	 0u                        C�	 ��                         ��	 <u                        ��	 ��                         :�	 Hu                        ��	 ��                         ��	 Tu                        '�	 ��        [                       ��	 `u                         
 ��                         P 
 lu                        � 
 Ȫ                         � 
 xu                        1
 Ъ                         x
 �u                        �
 ت                         
 �u                        M
 �                         �
 �u                        �
 �                         1
 �u                        }
 �                         �
 �u                        
 ��                         X
 �u                        �
 ��                         �
 �u                        1
 �                         y
 �u                        �
 �                         
 �u                        y
 �                         �
 �u                        1
 �                         �
 �u                        �
 �                \               !
 v                        q
  �                         �
 v                        	
 (�                         u	
  v                        �	
 ,�                         ^

 ,v                        �

 0    	                    
 0                          5
 �    	                    i
 �         �
                          �
           �
                         &
          Q
                          �
           �
 p    	                    �
 p         
 �    	                    C
 �         q
 `                        �
 `         �
 P
                         
 P
         +
 @
                        \
 @
         �
 �W                       �
 �W         �
 ��     h                   �
 �[                       '
 �[         K
 `�     h                   s
 �    	 ]                         �
 �         �
 �    	                    �
 �         
 @3                       ?
 @3         ]
 ��     H                   
 �L                        �
 �L         %
 �                        V
 �         �
 �                        �
 �         �
 P�    "                    �
 P�         �S               �R               
 `�	                       T
 `�	         �
 ��     0                   �
 ��	                       '
 ��	         j
  �     0                   �g               �
 �I	                       �
 �I	         9
  �     x                   ~
 �J	                       �
 �J	         
  �     `                   K
 `L                       q
 `L         �
 ��                         �
 �r	                       �
 �r	         ?
 ��     (                   �
 �q	            ^                 �
 �q	         
  �     P   	                U
  7                       �
  7         �
 �4                       ?
 �4         �S               2S               �
 �W    $                   �
 �W         �
 p[    $                   
 p[         %
 0�	    $                   n
 0�	         �
 P�	    $                   �
 P�	         �g               =
 3    $                   a
 3         
 �I	    $                   �
 �I	         
 �J	    $                   N
 �J	         �
 0L    $                   �
 0L         �
 �r	    $                   
 �r	         _
 `q	    $                   �
 `q	         �
 �6    $                   9
 �6         �
 �4    $                   �
 �4         
 p    #                   L
 p         u
 �	    #                   �
 �	         �
 �    #               _          �
 �         
 �    #                   I
 �         u
 p    #                   �
 p         �
 @    #                    
 @         9 
 0    #                   k 
 0         � 
 �    #                   � 
 �         � 
 �    #                   -!
 �         [!
     #                   �!
          �!
 @    #                   �!
 @         �!
 0i	    (                   "
 0i	         #"
 ��     8                   ="
  i	    0                   Y"
  i	         o"
 `H	    (                   �"
 `H	         �"
 `�     8                   �"
 0H	    0                   �"
 0H	         �"
 `+    (                   #
 `+         *#
 0+    0                   N#
 0+         l#
 �    (                   �#
 �         �#
 `    0                   �#
 `         �#
 �    T                   $
 �         &$
 `      ��                         D$
 Т                       d$
 Т         ~$
 �
                       �$
 �
         �$
  �     X   
                �$
 �
    $                   
%
 �
         )%
 �C         k%
 0�    �                  �%
 0�         �%
 ��    1  	                �%
 ��         ��              &
 @o    t                   F&
 @o         k&
 �n    t                   �&
 �n         �&
 Pp    ]                   �&
 Pp         '
 �v    t                   6'
 �v         ['
 v    t                   �'
 v         �'
 �w    ]                   �'
 �w         �'
 0�    L                   (
 0�         ;(
 ��     h                   \(
 @�    L                   (
 @�         �(
 ��    H                   �(
 ��         )
 ��    H                   Y)
 ��         �)
 ��    G                   �)
 ��         �)
 ��    a      G                   *
 ��         (*
 �    #                   Y*
 �         �*
 �    #                   �*
 �         �*
 �    N                   +
 �         0+
      N                   _+
           �+
 p    N                   �+
 p         �+
      N                   ,
           @,
 �    #                   o,
 �         �,
 �    #                   �,
 �         �,
 �    #                   -
 �         D-
  �    L                   g-
  �         �-
  �     h                   �-
 �    L                   �-
 �         �-
 `�    H                   &.
 `�         a.
 p�    H                   �.
 p�         �.
 ��    G                   /
 ��         '/
 ��    G                   O/
 ��         q/
 
    #                   �/
 
         �/
      #                   �/
           )0
 �    N    b                     T0
 �         y0
 `	    N                   �0
 `	         �0
 �
    N                   1
 �
         -1
 `
    N                   ^1
 `
         �1
 �	    #                   �1
 �	         �1
 0	    #                   2
 0	         72
  	    #                   e2
  	         �2
 �U    �                   �2
 �U         �2
  T    �                   3
  T         53
 �V    �                   c3
 �V         �3
  U    �                   �3
  U         �3
 �W                       4
 �W         /4
 �Y    �                   \4
 �Y         �4
 �W    �                   �4
 �W         �4
 �Z    �                   5
 �Z         -5
 �X    �                   [5
 �X         �5
 �[                       �5
 �[         �5
 �	                       6
 �	         ]6
 ��	                       �6
 ��	         �6
 p�  c        k                    Z7
 p�         �7
  �    k                    B8
  �         �8
 p�	                       9
 p�	         E9
 0�	                       �9
 0�	         �9
 �	                       :
 �	         ]:
 ��    ^                    �:
 ��         ;
 p�    S                    |;
 p�         �;
 ��	                       *<
 ��	         m<
 �A    X                   �<
 �A         �<
 pA    X                   �<
 pA         �<
 �B    R                   =
 �B         9=
 �o	    I                   U=
 �o	         k=
 ��     H                   �=
 �n	    I                   �=
 �n	         �=
  o	    E                   �=
  o	         >
 0n	    E                   M>
 0n	         {>
 po	    G                   �>
 po	         �>
 �n	    G                   �>
 �n	         �>
 p    #                   ?
 p         5?
 �    #   d                      _?
 �         �?
 �    N                   �?
 �         �?
 @    N                   �?
 @         @
 �    N                   ,@
 �         K@
 P1    �                   r@
 P1         �@
 �/    �                   �@
 �/         �@
 02    �                   A
 02         %A
 p0    �                   MA
 p0         oA
 P3                       �A
 P3         �A
 pI	                       �A
 pI	         9B
 PI	                       �B
 PI	         �B
 ��    _                    /C
 ��         �C
 ��    _                    D
 ��         mD
 ��    _                    �D
 ��         CE
 @�    _                    �E
 @�         F
  �    _                    �F
  �         �F
 �I	                       8G
 �I	         yG
 �J	                       �G
 �J	         H
 pJ	                       HH
 pJ	         �H
 � e         ;                    �H
 �         7I
     >                    �I
          �I
 P    M                    ?J
 P         �J
 �    <                    �J
 �         EK
 �J	                       �K
 �J	         �K
 p�    U                   �K
 p�         L
 �    U                   'L
 �         AL
 @�    Q                   zL
 @�         �L
 ��    Q                   �L
 ��         M
 ��    �                   >M
 ��         ]M
 �    �                   �M
 �         �M
 `                        �M
 `         N
 �                        4N
 �         aN
                          �N
           �N
 P                        �N
 P         )O
 �                        TO
 �         yO
 `    B                    �O
 `         �O
 �    Q                    �O
 �         /P
 �    �                    [P
 �       f        �P
      �                    �P
           �P
 P�    T                   Q
 P�         'Q
 0J    �                  MQ
 0J         mQ
 0H    �                  �Q
 0H         �Q
 pL                       �Q
 pL         �Q
 `r	                       AR
 `r	         �R
 @r	                       �R
 @r	         S
 P�    Z                    nS
 P�         �S
 �r	                       T
 �r	         ST
 p6                       �T
 p6         �T
  �     (                   AU
 6                       �U
 6         �U
 �6                       5V
 �6         �V
 P6                       �V
 P6         %W
 7                       uW
 7         �W
 @q	                       X
 @q	         IX
  q	                       �X
  q	         �X
  G    #                   &Y
  G         sY
  z    _                    �Y
  z         YZ
 �yg          _                    �Z
 �y         ?[
 0L    _                    �[
 0L         -\
 �L    _                    �\
 �L         ]
 �z    _                    �]
 �z         ^
 �q	                       M^
 �q	         �^
 p4                       �^
 p4         /_
 ��     P   	                }_
 04                       �_
 04         `
 �4                       q`
 �4         �`
 P4                       a
 P4         aa
 �4                       �a
 �4         �a
 �h	    B                   b
 �h	         -b
 h	    B                   Ib
 h	         _b
 `h	    B                   �b
 `h	         �b
 �g	    B                   �b
 �g	         �b
      #                   c
           -c
 P    #                   ^c
 P         �c
 �    ,                    �c
 �         d
 �                       "d
 �         =d
 `i	    h      (                   Yd
 `i	         od
 �                        �d
 �         e
 �    "                   3e
 �         _e
 p*    �   
                �e
 p*         �e
 P�     8                   �e
 �)    �   
                �e
 �)         f
  +                       9f
  +         [f
 `*                       �f
 `*         �f
 �+    (                   �f
 �+         �f
 ��         g
 ��         %g
 �    �                   Mg
 �         og
 �    �                   �g
 �         �g
 �	    �                   �g
 �	         h
      �                   .h
           Qh
 �
                       vh
 �
         �h
 �G	    B                   �h
 �G	         �h
 PG	    B                   �h
 PG	         �h
 �G	    6                   i
 �G	         )i
 G	    6                   Fi
 G	         ]i
 @�                        �i
 i      @�         �i
 ��                        �i
 ��         �i
 �    #                   !j
 �         ?j
 �H	    (                   Zj
 �H	         oj
 �    �                   �j
 �         �j
 ��     8                   �j
 �    �                   �j
 �         k
 �    �                   Ck
 �         dk
 �    �                   �k
 �         �k
 �    (                   �k
 �         �k
 ��	    V                   l
 ��	         Hl
 p    �                  �l
 p         m
  M    �                  �m
  M         n
 PJ    �                  |n
 PJ         �n
 ��	    V                   %o
 ��	         To
 P�	    V                   �o
 P�	         �o
 �#                         �o
 `~                        �o
 P�	    V                   p
 P�	         Jp
 �$                         fp
 �                        �p
 �=    j      �  "                �p
 �=         �p
 ��	    V                   Eq
 ��	         �q
 0$                         �q
 �~                        *r
 �	    V                   �r
 �	         �r
 $                         )s
 �~                        ns
 P�	    V                   �s
 P�	         �s
 @                         t
 Ps     8                   "t
 �p    Q  ,                ^t
 �p         �t
 �	    V                   �t
 �	         u
 0                         'u
 s     8                   Hu
 `i    Q  ,                �u
 `i         �u
 P�	    V                   v
 P�	         vv
 %                         �v
 ��                        w
 ��	    V                   gw
 ��	         �w
 �$                         x
 @�                        Rx
 �	    V                   �x
 �	         �x
 `                         �x
 �s         k                     �x
 ��    �                   ^y
 ��         �y
 ��	    V                   z
 ��	         vz
 �$                         �z
 ��                        {
 �	    V                   d{
 �	         �{
 �$                         |
 0�     8                   L|
 ��	    V                   �|
 ��	         �|
 p$                         �|
 p     8                   �|
 0�	    Q                   }
 0�	         :}
 �	    Q                   l}
 �	         �}
 ��	    Q                   �}
 ��	         �}
 ��	    Q                   #~
 ��	         N~
 0�	    Q                   �~
 0�	          
 p�	    Q                   \
 p�	         �
 ��	    Q                   �
 ��	         �
 ��	    Q                   z�
 ��	         Ҁ
 �	    Q                   0�
 �	         ��
 p�	    Q                   ��
 p�	         �
 0�	    Q            l             I�
 0�	         ��
 p�	    Q                   ��
 p�	         T�
 �	    Q                   ��
 �	         ��
 ��	    �                   �
 ��	         �
  �    �                   t�
  �         ҄
 ��    P                   =�
 ��         ��
 p�    �  +                �
 p�         ��
 ��    �  +                �
 ��         z�
 ��    �                  ڇ
 ��         4�
 0�    ^                   ��
 0�         
�
 �}    �                  M�
 �}         ��
      <                   �
           F�
 `�	    �                    ��
 `�	         ��
  �	    �                    �
  �	         *�
 �                      q�
 �         ��
 �                      ��
 �         �]              :�
 �    j                  ��
 �         �
 P
    6                   i�
 P
         ��
 �    [                   �
 �         m      n�
 �    �                  ˎ
 �         "�
 ��    �                  ��
 ��         �
 �
    6                   Q�
 �
         ��
      [                   �
           V�
 ��    j                  
 ��         (�
 �
    8                   ��
 �
         ܒ
 `    [                   6�
 `         ��
 ��                      ��
 ��         \�
     8                   ��
          �
 `    �                   o�
 `         ȕ
 �    [                   "�
 �         v�
 ��    �                  �
 ��         N�
 �	    H                   ��
 �	         �
 �     �                  q�
 �          ژ
 �	    Q                   7�
 �	         7^              ��
 �R    �                  �
 �R         ��
 0l    �                  �
 0l         ��
 �O    �                  �
 �O         ��
 `U    K         n               �
 `U         ��
 �X    |                  �
 �X         ��
 �H    �                  �
 �H         z�
 0G    �                  ��
 0G         h�
 �w    �                  ޠ
 �w         N�
 �u                      ��
 �u         .�
 ��    �  &                ��
 ��         "�
 �                      ��
 �         ��
 ��                      o�
 ��         ڤ
 ��                      K�
 ��         ��
 �    H	                  7�
 �         ��
 ��    [                   #�
 ��         ��
 ��    |                   ��
 ��         d�
 ��                      ը
 ��         @�
 0�    �                  ��
 0�         <�
 P�    [                   ��
 P�         �
 ��    |                   ��
 ��         �
 @�    �                  o�
 @�         �
 0�    [                   [�
 0�         ƭ
  �    | o                        4�
  �         ��
 `�    �                  �
 `�         ��
 ��    [                   	�
 ��         t�
  �    |                   �
  �         J�
  �    �	                  ˱
  �         F�
 ��    [                   ��
 ��         "�
  �    |                   ��
  �         ��
 ��    �                  y�
 ��         ��
 �    [                   e�
 �         е
  �    �                   B�
  �         ��
 ��    |                   �
 ��         ��
 ��    2  %                �
 ��         ��
 ��    2  %                �
 ��         ��
 �    �                  ��
 �         b�
 �    �  	                �
 �         \�
 �o    �  	                ӻ
 �o         D�
 0�	         r�
 �                         ��
                           ��
                           �
 @                         R�
 �p                               p�
 `                         ��
 �                         �
                           $�
                           n�
 �                         ��
 �                         ־
 @                         �
 ��                         �
 ��                         -�
 Pw                        N�
 �                         h�
 ��                         ��
 x                        ��
 �     :                    �
 `�     :                    6�
 ��                         Z�
 Py                        ~�
 ��                         ��
 ��                         ��
 `�                         ��
 У                         ��
 @�                         �
 w                        >�
 @�                         f�
 �y                        ��
 `�                         ��
 �y                        ��
  �     q      <                    %�
 ��     <                    l�
 ��     ;                    ��
 ��     C                     �
 �x                        N�
 @�     ;                    ��
  �     C                    ��
 Px                        0�
 `�                         R�
 �w                        t�
 ��     �                   ��
 @�     X                   ��
 �W                         ��
 �W                         "�
 �W                         H�
 pW                     .text   �                       .data                           .bss    P                            n�
 0�                         ��
 8v                        ��
 4�                         �
 Dv                        B�
 8�                         u�
 Pv                        ��
 <�                         ��
 \v                        �
 @�                         >�
 hv           r                   p�
 D�                         ��
 tv                        ��
 H�                         �
 �v                        D�
 L�                         w�
 �v                        ��
 P�                         ��
 �v                        �
 T�                         @�
 �v                        r�
 X�                         ��
 �v                        ��
 \�                         ��
 �v                        �
 `�                         L�
 �v                        z�
 d�                         ��
 �v                        ��
 h�                         ��
 �v                         �
 l�                         w�
 �v                        ��
 p�                          �
 �v                        2�
 t�                         W�
 w                        |�
 x�                         ��
 w                  s            ��
 |�                         �
 w                        `�
 ��                         ��
 (w                        ��
 ��                         <�
 4w                        ��
 ��                         ��
 @w                        �
 ��                         ;�
 Lw                        b�
 ��                         ��
 Xw                        ��
 ��                         =�
 dw                        ��
 ��                         ��
 pw                        (�
 ��                         y�
 |w                        ��
 ��                         ��
 �w                         �
 ��                         K�
 �w                        v�
 ��                         ��
 �w                        
�
 ��                         T�
 �w                        ��
 ��                         ��
 �w                        ��t      
 ȫ                         0�
 �w                        x�
 Ы                         ��
 �w                        �
 ث                         /�
 �w                        V�
 �                         ��
 �w                        ��
 �                         1�
 �w                        z�
 �                         ��
  x                        �
 ��                         m�
 x                        ��
  �                         ��
 x                        �
 �                         N�
 $x                        ~�
 �                         ��
 0x                        ��
 �                         �
 <x                        6�
  �                         k�
 Hx                        ��
 (�                         ��
 Tx                        
�
 0�                         =�
 `x                        p�
 8�   u                            ��
 lx                        ��
 @�                         �
 xx                        D�
 H�                         m�
 �x                        ��
 P�                         ��
 �x                        ��
 X�                        �
 �x                        $�
 h�                        A�
 �x                        ^�
 x�                        z�
 �x                        ��
 ��                        ��
 �x                        ��
 ��                        ��
 �x                        �
 ��                        =�
 �x                        b�
 ��                        ��
 �x                        ��
 Ȭ                        ��
 �x                        ��
 ج                        �
 �x                        4�
 �                         U�
 y                        v�
 ��        v                       ��
 y                        ��
 ��                         ��
  y                        �
 �C    H                     V�
  �                          ��
 ,y                         ��
 �     `                   �
 8y                        D�
 h�     .                   v�
 Dy                    .rdata        �  M                 ��
 ��                         ��
 Py                         �
 ��                         ,�
 \y                        X�
 ��                         ��
 hy                        ��
 ��                         ��
 ty                        �
 ��                         4�
 �y                        `�
 ��                         ��
 �y                        ��
 ��                        ��
 �y                         �
 ԭ                        $�
 �y                        H�
 �               w               ��
 �y                        ��
 �                        �
 �y                        P�
 (�                        y�
 �y                        ��
 D�                        ��
 �y                        ��
 `�                         &�
 �y                        X�
 d�                         ��
 �y                        ��
 h�                         ��
 �y                        �
 p�                         D�
 z                        t�
 x�                         ��
 z                        ��
 ��                         
�
 z                        <�
 ��                         l�
 (z                        ��
 ��                         ��
 4z                        ��
 ��                         )�
 @z                        X�
 ��                        |�
 Lz                        ��
 ��                      x        ��
 Xz                        ��
 ̮                        *�
 dz                        l�
 �                        ��
 pz                        ��
 �                        �
 |z                        B�
  �                        k�
 �z                        ��
 <�                         ��
 �z                        ��
 @�                         *�
 �z                        \�
 D�                         ��
 �z                        ��
 L�                         ��
 �z                        �
 T�                         F�
 �z                        x�
 \�                         ��
 �z                        ��
 d�                         �
 �z                        <�
 h�                         k�
 �z                        ��
 l�                         ��
 �z                        ��
 p�     (                   &�
  {y                              T�
 ��     (                   ��
 {                        ��
 ��     (                   ��
 {                        �
 �     (                   =�
 ${                        l�
 �                         ��
 0{                        ��
 �     (                   ��
 <{                        �
 <�     (                   L�
 H{                        z�
 d�     (                   ��
 T{                        ��
 ��     (                   �
 `{                        6�
 ��                         a�
 l{                        ��
 ��                         ��
 x{                         �
 ��                         j�
 �{                        ��
 ��                         &�
 �{                        ��
 Ȱ                         �
 �{                        ��
 а                         ��
 �{     z                         (�
 ԰                         r�
 �{                        ��
 ذ                         �
 �{                        P�
 ܰ                         ��
 �{                        �
 �                         x�
 �{                        ��
 �                         .�
 �{                        x�
 �                         ��
 �{                        ��
 ��                         ��
 �{                        �
 ��                         6�
 |                        \�
  �                        y�
 |                        ��
 �                        ��
  |                        ��
 8�                        �
 ,|                        :�
 T�                        o�
 8|                        ��
 p�                        ��
 D|                        ��
 ��                        �
 P|           {                    �
 ��                         K�
 \|                        v�
 ��                         ��
 h|                        ��
 ��                         ��
 t|                        �
 ��                         ;�
 �|                        `�
 ��                         ��
 �|                        ��
 ȱ     (                   ��
 �|                        ��
 �     (                   $�
 �|                        L�
 �     (                   u�
 �|                        ��
 @�     (                   ��
 �|                        ��
 h�                         �
 �|                        :�
 l�                         ��
 �|                        ��
 p�                         �
 �|                        Z�
 t�                         ��
 �|                        8  |�                         �  �|                  |             ��                         � }                        � ��                         c }                        � ��                         B }                        � ��                         � (}                        B ��                         � 4}                        � ��                          @}                        b ��                         � L}                         ��                         s X}                        � ��                         ) d}                        � ��                         � p}                        > Ȳ                         � |}                        � ̲                        � �}                        	 �                        1	 �}                        R	 �                        �	 �}                        �	}        �                         
 �}                        :
 <�     4                   `
 �}                        �
 p�     4                   �
 �}                        �
 ��                          �}                        : ��                         n �}                        � ��                         � �}                         ��                         G �}                        z ��                         �  ~                        � ��                         � ~                        ( ��                         ` ~                        � ��                         � $~                        � ĳ                         , 0~                        f ȳ                        � <~                        � ܳ                         � H~                        � �   ~                             T~                        D �                         k `~                        � �                         � l~                        $ �                         m x~                        � �                          �~                        z ��                         � �~                         ��                         ` �~                        �  �                          �~                        \ �                         � �~                         �                         [ �~                        � �                          �~                        R �                         � �~                        � �                         - �~                        v �                         � �~                         �                               � �~                         $�                         �                         � ,�                         u                         � 4�                         m                          � <�                         a ,                        � D�                         ! 8                        j H�                         � D                         L�                         f P                        � P�                          \                        d T�                         � h                         X�                         _ t                        � \�                        � �                        � x�                          �                        $  ��                        F  �                        h  ��               �               �  �                        �  ̴                         �  �                        
! д                         <! �                        n! Դ                         �! �                        �! ܴ                         " �                        2" �                        O" �                        l" �                         �" �                        # ��                         9# �                        l# ��     &                   �# �                        �# $�     &                   �# �                        $ L�                         5$ �                        ^$ P�                         �$ (�                        �$ T�                        �$ 4�                        �$ ��                        % d�                          E% @�                       �        k% h�     &                   �% L�                        �% ��     &                   �% X�                        & ��     &                   9& d�                        c& �     &                   �& p�                        �& �                         �& |�                        ' �                        ' ��                        ;' (�                        W' ��                        s' D�                         �' ��                        �' L�                         �' ��                        �' T�                         ( ��                        G( X�                         q( Ā                        �( `�                         �( Ѐ                        �( d�                        ) ܀                        ) t�     (                   D) �                        k) ���           (                   �) �                        �) Ķ     (                   �)  �                        	* �     (                   1* �                        Y* �                        }* �                        �* $�                         �* $�                        + ,�                         k+ 0�                        �+ D�                         P, <�                        �, \�                         J- H�                        �- t�                         �- T�                        1. |�                         e. `�                        �. ��                         �. l�                        / ��     �                   :/ x�                        q/ �                         �/ ��                        10  �                         �0 ��                        �0 (�     �                          -1 ��                        i1 0�     �                   �1 ��                        �1 �                         2 ��                        [2 ��     �                   �2 ��                        �2 ��                         73 ́                        �3 ��                         �3 ؁                        ]4 ȹ                         �4 �                        �4 й                         45 ��                        �5 �                         �5 ��                        [6 �                         �6 �                        7 ��                         R7 �                        �7  �                         �7  �                        �7 �                         8 ,�                        K8 �                         |8 8�                        �8 �            �                   �8 D�                        9  �                         n9 P�                        �9 (�                         (: \�                        �: 0�                         �: h�                        �: 8�                         V; t�                        �; @�                         < ��                        s< H�                         �< ��                        �< P�                         == ��                        �= X�                         �= ��                        W> `�                         �> ��                        �> h�                         �> ��                        #? x�                         �? Ȃ                        �? ��                         Y@ Ԃ                        �@ ��     |                   ?A ��                        �A �     |             �            3B �                        �B ��     9                   C ��                        oC Ȼ                         �C �                        MD л                         �D �                        �D �                         7E �                        �E �                         �E (�                        F ��                         PF 4�                        �F  �     <                   �F @�                        G <�     <                   eG L�                        �G x�                         H X�                        �H ��                         �H d�                        CI ��                         �I p�                        �I ��                         WJ |�                        �J ��                         "K ��                        �K Լ                         �K�       ��                        KL ܼ                         �L ��                        M �                         nM ��                        �M ��                         9N ��                        �N �                         �N ă                        MO �                         �O Ѓ                        'P $�                         �P ܃                        �P ,�                         CQ �                        �Q <�                         �Q �                        YR D�                          �R  �                        9S d�                         �S �                        �S l�                         eT �                        �T ��                         3U $�                        �U ��                         V 0�                        �V ��                          W <�   �                           �W ��                         )X H�                        �X ؽ                         'Y T�                        �Y �                         /Z `�                        �Z �                         2[ l�                        �[  �                         (\ x�                        �\ 8�                         ] ��                        �] P�                         ^ ��                        y^ l�     <                   �^ ��                        u_ ��     /                   �_ ��                        Y` ؾ     /                   �` ��                        =a �     /                   �a ��                        !b 8�     >                   �b ̄                        %c x�                         �c ؄                        	d ��                         xd �        �                      �d ��                         Ye ��                        �e ��     >                   Mf ��                        �f �                         Ag �                        �g �                         "h �                        �h �     >                   i  �                        �i 0�                         j ,�                        yj 8�                         �j 8�                        Wk @�     >                   �k D�                        [l ��                         �l P�                        ?m ��                         �m \�                        n ��     >                   �n h�                        !o ��                         �o t�                        p ��                         tp ��                        �p ��     >                   eq ��               �               �q  �                         Yr ��                        �r (�                         >s ��                        �s 8�                          t ��                        �t @�     6                   u ��                        �u x�     6                   v ȅ                        �v ��     0                   w ԅ                        �w ��     8                   x ��                        �x �                         �x �                        wy 0�	    �                    �y 0�                          �y ��                     .ctors  P�	                        -z ��                        tz ��                          �z �	                        �z �	         ?{ К                        �{ К         �{ P�                        | P�         [| 0�                        �| 0�       �        �|  �                        <}  �         �} `�                        �} `�         ~ @�                        a~ @�         �~ p	    a                   �~ p	         5 ��                        ��         � ��                       � ��         Q� P�    u                   �� P�         � ��    	                   8� ��         �� ��                        Ձ ��         �  �                        p�  �         �� �    (                   � �         K� Г    (                   �� Г         �  �                        6�  �         y�  �                        Ǆ  �         � ��    '                   Z� ��         �� ��    '                   � ��         /� 0	    %                    z� 0	         �� ��    '                   7� ��         �� p�    '                   !� p�               ��  �    '                   �  �         5� ��    '                   �� ��         ׉ ��                        "� ��         g� � 	    �                   �� � 	         �� �	    <                  F� �	         �� ��    i                   Ջ ��         � p		                        W� p		         �� p	                        ь p	         �  	                        O�  	         ��  	                        э  	         � �		                       U� �		         �� �	                       ێ �	         � �	    K                    ^� �	         �� �	    K                    ޏ �	         �  	    b                    c�  	         ��  	    b                    �  	         /� �		                       o� �		         �� �		                       � �		         #� �
	                   �          g� �
	         �� 
	    �                   � 
	         %� @�                        i� @�         �� И                        � И         +�  �                        m�  �         �� ��                        � ��         )� 0�                        n� 0�         �� P�                        � P�         3�  �    
                    v�  �         �� ��    
                    �� ��         5� 0�                        {� 0�         �� ��                        �� ��         =� П                        �� П         Ř �    
                    
� �         I� ��                        �� ��         ˙ @�                        � @�         Q� P�                        �� P�         ۚ 0�                        #� 0�         e� ��                      �� ��         � 0�    I      �                   8� 0�         � P�                        Ü P�         �  �    	                    F�  �         �� `�                        Ɲ `�         � `	                        A� `	         {� p�    &                   �� p�         �� ��    &                   :� ��         u�  �                        ��  �         �� �                        <� �         {� �                        �� �         �� ��                        ?� ��         }� 	    k                   �� 	         �� `	    h                   ?� `	         �� P�                       ʢ P�         � `�    �                   U� `�         �� ��    a                   ܣ ��         � p�    -                   �� p�         � ��    S                   V� ��         ��   	                       �   	         E� ��    �      .                  �� ��         � 0�    !                   '� 0�         g� `�    A                   �� `�         � P�                       2� P�         q� ��                        �� ��         �� 0	    )                   7� 0	         q� ��    @                   �� ��         ��  �    9                   e�  �         ˪ 0�    H                   � 0�         W� p�                       ȫ p�         3� @�    6                   �� @�         � �    �                  V� �         �� p�    M                   � p�         /� 0�                       w� 0�         ��  	    (                   �  	         _� ��                        �� ��         � ��    1                   V� ��         �� �    =                   � �         '� �
	    1                   i� �
	         ���       ��    @                   � ��         3� ��    <                   |� ��         �� P�    J                   � P�         Q�  �    \                   ų  �         3� P�    O                   �� P�         � ��    �                   a� ��         ��  �    s                   ��  �         ;� ��    b                   �� ��         � ��    b                   �� ��         � �    _                   �� �         � ��    G                   �� ��         �  �    b                   ��  �         �� ��    b                   n� ��         ݻ @�    V                   %� @�         g� ��    h                   �� ��         �� `�    w                   g� `�         ӽ   	    �                   �   	         c� ��                       �� ��         � �	                       3� �	  �             q� ��    D                   �� ��         � `�    -                   I� `�         �� �    H                   �� �         � p	    H                   U� p	         �� �	    7                   �� �	         7� ��    7                   �� ��         �� Ж    o                   .� Ж         o� 0�                       �� 0�         �� ��                        :� ��         y� @�                        �� @�         �� ��                        I� ��         �� ��    �                    �� ��         � P�                       d� P�         �� P�    0                   �� P�         /� `�    J                    t� `�         �� P�    �                    �� P�         ?� ��                       �� ��         ��  �    0                   �  �         W� �    1                    �      �� �         �� �    S                    0� �         }� ��    S                    �� ��         � @�    k                   l� @�         �� p�    J                    � p�         O� ��    S                    �� ��         �� ��                       =� ��         �� P�    0                   �� P�         #� �    1                    q� �         �� ��    ^                    � ��         a� `�    Y                    �� `�         � ��    y                   \� ��         ��  �    D                    ��  �         K� @�    N                    �� @�         �� ��                       E� ��         �� �    0                   �� �         7� ��    1                    �� ��         �� ��    �                     � ��         e� �    �                   �� �         �� ��             �               H� ��         �� ��    �                   �� ��         � 0�    �                   h� 0�         ��  �    �                   ��  �         ?� @�                        �� @�         ��  �                        5�  �         �� 0�                        �� 0�         #� �                        v� �         �� ��	    �                   � ��	         g� ��	    �                   �� ��	         � `�    �                   �� `�         #� �		                       �� �		         � �	                       s� �	         �� ��    �                   q� ��         �� @	                       F� @	         �� @	                       �� @	         � ��    �                   �� ��         ��  	                       -�  	         k�  	                       ��  	         �� ��	    ] �                        @� ��	         �� �		                       �� �		         #� �	                       q� �	         �� ��    �                   '� ��         �� `	    E                   �� `	         � `	    E                   g� `	         �� �	    L                   �� �	         1� �	    L                   w� �	         ��  		    L                   �  		         G�  	    L                   ��  	         �� �	                       � �	         a� �	                       �� �	         �� �	    A                   2� �	         s� �	    A                   �� �	         �� P		                       V� P		         �� P	                       � P	         [� �		                       �� �		         �� �	                       B� �	         �� p�    X                   �� p�         � �֔          
                    �� ��         �� ��    
                    g� ��         �� �[                     .text   �                       .data                           .bss    P                            � 4�                         `� �                        �� 8�                         �� �                        :� <�                         �� �                        �� @�                         � (�                        f� D�                         �� 4�                        � H�                         P� @�                        �� L�                         �� L�                        8� P�                         �� X�                    .rdata  �     �                    �� T�                         � d�                        h� \�                         �� p�                        �� `�     �                          I� |�                        �� d�                         �� ��                        0� p�                         �� ��                        �� t�                         )� ��                        z� x�                         �� ��                        � |�                         j� ��                        �� ��                         � Ć                        `� ��                         �� І                        �� ��                         C� ܆                        �� ��                         �� �                        *� ��                         v� �                        �� ��                         �  �                        Z� ��                         �� �                        L� ��                         �� �                        >� ��            �                   �� $�                        �� ��                         =� 0�                        �� ��                         �� <�                        *  ��                         w  H�                        �  ��                          T�                        ` ��                         � `�                        � ��                         3 l�                        t ��                         � x�                        � ��                         ; ��                        � ��                         � ��                        
 ��                         Q ��                        � ��                         � ��                        &  �                         j ��                        � �                         � ��                        6 �                   �             ̇                        � �                          ؇                        Z �                         � �                        � �                          ��                        ^ �                         � ��                        �  �                        ,	 �                        p	 0�                         �	 �                        �	 4�                         @
  �                        �
 8�                         �
 ,�                         <�                         P 8�                        � @�                         � D�                          D�                         g P�                        � H�                         � \�                        6 L�                         { h�                        � P�                         �       t�                        N T�                         � ��                        � X�                           ��                        h \�                         � ��                        � `�                         9 ��                        ~ d�                         � ��                         h�                         U ��                        � l�                         � Ȉ                        0 p�                         w Ԉ                        � ��                         ��                        Z ��                         � �                        � ��                         * ��                        p ��                         � �                        � ��                         5 �                        v ��                         � �   �                           � ��                         > (�                        � ��                         � 4�                        
 ��                         P @�                        � ��                         � L�                         ��                         c X�                        � ��                         � d�                        * ��                         s p�                        � ��                          |�                        P ��                        � ��                        � �                         ( ��                        n �                         � ��                        D �                         � ��                          $�                         h ��                        � (�                          ĉ        �                      T <�                         � Љ                        � D�                         ) ܉                        p L�                         � �                        � P�                         C  �                        �  X�                         �   �                        ! `�                         T! �                        �! h�                         	" �                        v" t�                         �" $�                        
# |�                         |# 0�                        �# ��                         \$ <�                        �$ ��                         % H�                        j% ��                         �% T�                        & ��                         K& `�                        �& ��                         �& l�               �               B' ��                         �' x�                        �' ��                         B( ��                        �( ��                         �( ��                        ") ��                         e) ��                        �) ��                         �) ��                        >* ��                         �* ��                        �* ��                         + ��                        l+ ��                         �+ ̊                        V, �                         �, ؊                        >- �                         �- �                        �- �                         ). ��                        v.  �                         �. ��                        `/ (�                         �/ �                        L0 0�                         �0 �                      �        Z1 8�                         �1  �                        ^2 @�                         �2 ,�                        \3 H�                         �3 8�                        H4 P�                         �4 D�                        �4 \�                         %5 P�                        p5 l�                         �5 \�                        V6 |�                         �6 h�                        �6 ��                         87 t�                        �7 ��                         �7 ��                        8 ��                         X8 ��                        �8 ��                         �8 ��                        69 ��                         ~9 ��                        �9 ��                         	: ��                        L: ��                         �: ��                        �: �ŝ                               V; ȋ                        �; ��                         �; ԋ                        B< ��                         �< ��                        �< ��                         = �                        \= ��                         �= ��                        �= ��                         5> �                        �> ��                         �> �                        ? ��                         `? �                        �? ��                         �? (�                        :@ ��                         �@ 4�                        �@  �                         A @�                        ZA �                         �A L�                        �A �                         9B X�                        �B �                         �B d�                        C �     �                          dC p�                        �C  �                         D |�                        ^D (�                         �D ��                        E 4�                         RE ��                        �E 8�                         �E ��                        FF <�                         �F ��                        �F @�                         =G ��                        �G L�                         �G Č                        ,H P�                         �H Ќ                        �H X�                         3I ܌                        �I `�                         �I �                        6J l�                         �J �                        �J p�                         4K  �                        �K t�                         �K �                        8L x�            �                   �L �                        �L ��                         5M $�                        �M ��                         �M 0�                         N ��                         nN <�                        �N ��                         O H�                        \O ��                         �O T�                        �O ��                         <P `�                        �P ��                         �P l�                        "Q ��                         wQ x�                        �Q ��                         !R ��                        vR ��                         �R ��                        S ��                         rS ��                        �S ��     "                   T ��                        rT ��                         �T ��                        U �                   �            �U ��                        >V  �                         �V ̍                        $W $�                         �W ؍                        
X (�                         �X �                        0Y 4�                         zY ��                        �Y 8�                         Z ��                        XZ <�                         �Z �                        4[ H�                         y[ �                        �[ L�                         \  �                        H\ P�                         �\ ,�                        �\ p�                         ?] 8�                        �] t�                         �] D�                        ,^ x�                         �^ P�                        
_ ��                         U_ \�                        �_ ��                         �_�       h�                        6` ��                         }` t�                        �` ��                         a ��                        Ra ��                         �a ��                        �a ��                         6b ��                        �b ��                         �b ��                        c ��                         ]c ��                        �c ��                         �c ��                        6d ��                         ~d Ȏ                        �d ��                         "e Ԏ                        ~e ��                         �e ��                        6f ��                         �f �                        �f ��                         &g ��                        vg ��                         �g �                        h ��                         zh �   �                           �h ��                         ci �                        �i ��                          �i  s	         j ��     (                   j  s	         0j �r	     .text   �                       .data                           .bss    P                        .rdata  �                          Dj ��                        bj ��                          �j (�                         �j  s	                        �j ��                          �j 4�                         �j �r	    )                    
k ��                          %k @�                         @k P                          Wk 0K	         jk `�     (                   �k 0K	         �k  K	     .text   �                       .data                           .bss    P                        .rdata  �                          �k P                        �k ��        �                        �k L�                          l 0K	                        l  �                          3l X�                         Ml  K	    )                    fl �                          �l d�                         �l ��                          �l ��         �l ��     (                   �l ��         �l `�     .text   �                       .data                           .bss    P                        .rdata  �                          m ��                        0m �                          Qm p�                         rm ��                        �m �                          �m |�                         �m `�    )                    �m �                          n ��                         n ��                          Xn `�         �n 0�         �n �     X   
                �n 0�         o  �         Ao �� �              �o P�         �o  �         @p Ц                         Xp ��                        pp ��     "                    �p �b                    .text   �                       .data                           .bss    P                            �p ��    X                     
q �                          Kq ��                         �q `�                         �q $�                          'r ��                         ur 0�                        �r (�                          �r ��                         �r  �    )                    +s ,�                          Ys ��                         �s ��    v                    �s 4�                          jt ď                         �t P�    .                    3u D�                          �u Џ                         �u  �    I                    ,v P�                        �        vv ܏                     _ZdlPv  ��	                      .text   �                       .data                           .bss    P                            �v ��	                        �v `�                          �v �                     _ZdlPvy ��	                      .text   �                       .data                           .bss    P                            �v ��	                        �v d�                          w �                     _ZdaPv  ��	                      .text   �                       .data                           .bss    P                            w ��	                        "w h�                          0w  �                         >w ��	                      .text   �                       .data                           .bss    P                            Mw ��	                        bw l�                          xw ��                               �                                /               C               3               �               �           __tcf_0 ��	         �w @          �%               �w �         �w P�         
x P�         $x ��	         9x ��	         \x ��	         {x  �	         �x  �	     .text   �                       .data                           .bss    P                        .rdata  �     N                     �  ��	                        �  |�                         	  �                         �x �    Z                   �x ��     %                     y $�                         Ry P�                       �y ��     %                    �y 0�                         �y P�    %                    z ��                          1z <�                         Rz  �	    V                    qz ��                         �z H�     �                          �z ��	    )                    �z ��                         �z T�                         { ��	    H                    -{  �                         W{ `�                         �{ ��	    %                    �{ �                         �{ l�                         �{  �	    q   
                 )| �                          a| x�                     .ctors  X�	                        �| @                           �| `�	                          �| ��	         �| `�	         } 0R                        /} `{                        S} ��                         w} @K                    .text   �                       .data                           .bss    P                            �} `�	    3                    �} $�                          �} ��                         �} ��	    3                    �} ,�            �                    ~ ��                         .~ `�	    3                    U~ 4�                          }~ ��                         �~ ��	                          �~ ��	         �~  �	         �~ ��	         �~ ��	     .text   �                       .data                           .bss    P                             ��	                         2 <�                          Q ��                         p ��	    }                    � @�                          � ��                         �  �	    ~                    � H�                          � ��                         � ��	                        � P�                          ?� ̐                         `� ��	                        �� X�                          �� ؐ                         ŀ P�	                          ـ P�	         � �         � �         � P�    �           7� P�         R� �:         o� �:         �� @�	         �� p         �� �         � �         � �         +� P�         T� P�         }� @�         �� �         ��  �         ۂ  �     $                    
� c                        9� @�     (                   Q� ��     (                   n� ��     (                   �� P�     (               .text   �                       .data                           .bss    P                            ȃ P�	                         � `�                          �� �                         � �                         7� d�                          W� �                     .rdata        "                     w� P�                        �� h�                          �� ��                         ӄ �:                        �� l�                          � �         �                      >� @�	    
                    X� p�                          s� �                         �� p    
                    �� t�                          ͅ  �                         � �                         � x�                          D� ,�                         p� �    
                    �� |�                          ǆ 8�                         � P�                         "� ��                          R� D�                         �� @�    
                    �� ��                          � P�                         � �                         /� ��                          N� \�                         m�  �                         �� ��                          �� h�                         ؈ ��	                          � �.          �  �	     .text   �                       .data                       �          .bss    P                            5� ��	                        M� ��                          f� t�                         �  �	                        �� ��                          �� ��                         ؉ �.                           � ��                          <� ��         j� 0�         �� �         Ҋ  �         ��  �         9� �         �� ��	         �� ��	     .text   �                       .data                           .bss    P                            �� ��    ]                     � ��                          � ��                         J� ��    b                    ~� ��                          �� ��                         � 0�    S                   � ��                      .rdata  0     4                    G� ��                         w� �    �                    �� ��                          �      � ��                         H�  �    �                    w� ��                          �� ��                         ׎  �    �                    � ��                          `� ȑ                         �� �    �                   �� ��     8                    V� ԑ                         �� ��	    �                    ː �     4                    � ��                         � ��	                        "� L�                          @� �                         ^� ��                          �� �	         �� �H                        Ƒ а         � ��	         ��  I                        2� �	         K�  �	         `� ��	         z� p�	     .text   �                       .data                           .bss    P                            �� ��    9                    �� T�     -                    � ��               �                � �	                        #� ��                          :� �                         Q� а                        {� ��                          �� �                         ѓ ��	                        � ��                          � �                         � �	                        :� ��                          Z� (�                         z�  �	                        �� ��                          �� 4�                         ͔ ��	                        � ��                          � @�                         /� p�	                        K� ��                          h� L�                     .text   �                       .data                           .bss    P                            �� �                         �� �                          ��  �	         � ��	          � ��	     .text   �       �                      .data                           .bss    P                            .� �    @                    z� ��                          ǖ X�                         �  �	    X                    7� ��                          [� d�                         � ��	    s                    �� ��                          �� p�                         �� ��	    O                    ˗ ��                          �� |�                     .text   �                       .data                           .bss    P                            �� �                         �                                /               "� ��                       ]� ��         �� ��                       Ș ��         �� p�         � �          1� �          S� P�         z� @          �� �          C               �� 0�                       � 0�         � `��           (                   3               H� ��                       � ��         �� ��     (                   �               �  �    )                   �  �         �               E� ��    )                   |� ��         �� ��	         �%               ٛ  �    /                   �  �         I� �d                        �� ��	         �� @.          ��  .          � `d                        � �	         1� 0�	         E� `�     ,                    |� ��     '                .text   �                       .data                           .bss    P                        .rdata  p     �                     �� ��                         � ��                        &� ��                         ]� ��                        �� p�                        �� ��                          ՞ ��                         �� P�    �                          #� ��                          Q� ��                         � ��                         �� ��                        � ��                         � Ē                        U� ��                         �� В                        �� ��                         � ܒ                        +� ��	    D                    f� ��                         �� �                         ޡ �                         � ��                        V� ��	    P                   p� �     0                    ��  �                         �� �	    �                    �� @�     5                    ע �                         � 0�	    �                    
� x�     5                    %� �                         @�  .                          r� @                          �� �                          �� @.            �                    � �                          � �                          <� ��	                          W� `          y� ��	     .text   �                       .data                           .bss    P                            �� ��	                        �� ��                          Ӥ $�                         �� ��	                        � ��                          0� 0�                         N� `                          v� ^                      _Znwy   ��	                      .text   �                       .data                           .bss    P                            �� ��	    m                    �� ��                          �� <�                     _Znay   ��	                      .text   �                       .data                           .bss    P                            �� ��	                        �� ��                    �            ɥ H�                         ֥ ��	                      .text   �                       .data                           .bss    P                            � ��	                        � ��                          � T�                         :� `�	                          M� ��	     .text   �                       .data                           .bss    P                        .rdata        ?                     c� `�	    !                    |� ��                          �� `�                         �� ��	    !                    ̦ ��                          � l�                         � ��                          0� ��     X   
                `� ��         �� `�         �� ��         � ��         �� p�         �� `�     %                    *�  c                    .text   �                       .data                           .bss  �        P                            Z� ��                        �� ��                          �� x�                         � `�    )                    � ��                          M� ��                         ~� ��    a                    � ��                          G� ��                         �� ��    �                    2� ��                          �� ��                         @� p�    I                    �� �                          � ��                         �� ��	                          �� ��	         �� p�         ׮ p�         �� `�         @� ��	         T� ��         l� P�         �� 0�     @               .text   �                       .data                           .bss    P                            �� ��	                         į �                          ߯ ��                         �� p�                 �              #� �                          M� ��                         w� `�                         °  �                          � ̓                         Z� ��	    
                    t� $�                          �� ؓ                         �� ��    7                    ȱ (�                          � �                         � P�                        2� 0�                          _� �                         �� б                          �� �     X   
                � б         � ��         >� ��         �� 0�         � P�         �� ��     &                    �� @c                    .text   �                       .data                           .bss    P                            � б                        � 4�                          L� ��                         ~� ��    )                    �� 8�        �                        � �                         � ��    �                    x� @�                          ޶ �                         D� 0�                       �� T�                          #�  �                         �� P�    y                   � l�                          �� ,�                         *� ��                          W� p.      .text   �                       .data                           .bss    P                        .rdata  `     �                     �� ��    �                   ƺ ��     <                    �� 8�                         .� p.                          } �                         p� `�                          �� ��         �� д         ޻ д         �� �         5� ��         h� ��         �� �         �� @�         ؼ p�         �� �         � �         0� �         K� @� �              m� ��         ��  �         �� в         � б         � `�     .text   �                       .data                           .bss    P                        .rdata          =                 +� `�    �                    b� ��                          �� D�                         Ҿ ��    V                    �� ��                          � P�                         F� д                         i� ��                          �� \�                         �� �    o                    � ��                          2� h�                         s� ��    s                    �� ��     !                    �� t�                          � ��    P                    X� �                          �� ��                         �� �                         �� �                          � ��                         D� @�    & �                         f� �                         �� ��                         �� p�                         �� 8�                          �� ��                         � �    X                    ?� <�                          e� ��                         �� �                        �� D�                          �� ��                         �� @�    T                    � H�                          A� Ȕ                         j� ��    $                    �� X�                          �� Ԕ                         ��  �    \                    � d�                          F� ��                         v� в    :                    �� t�     !                    �� �                         � б                        A� ��                          f� ��                         �� `�    i                    �� ��              �                  �� �                         � `�	                          <� 0�	         p� @�	         ��  �         �� ��         � �         +� ��         Z� �U      .text   �                       .data                           .bss    P                        .rdata        �                     z� `�	                       �� ��     -                    �� �                         *� 0�	                       d� ��     -                    �� �                         �� @�	                       � �     -                    O� (�                         ��  �    ;                    �� 8�                          �� 4�                         1� ��                         c� D�                          �� @�                         �� �                         �� H�                          *� L�                         [� ��    �                           �� L�                          �� X�                         �� X                          � �U     0                    G� ��                          x� ��         �� `�         �� `�          � p�         #� p�         H� ��         p� ��         ��  �         �� �C	         �� `�     X   
                �� PR                        &� �C	         =�  E	         T� ��     X   
                o� `R                        ��  E	         �� �C	         �� �D	         �� `C	         �� `C	         �  C	         /�  C	         H� �D	         _� �D	         v� @D	         �� @D	     .text   �                       .data                           .bss    P                            �� ��                         �� P�                          � d�                         O� `�                         �� T�            �                    �� p�                         �� p�                         � X�                          :� |�                         d� ��                         �� \�                          �� ��                         �� ��                         � `�                          M� ��                         |�  �                         �� d�                          �� ��                         � �C	    Z                    %� h�                          C� ��                         a�  E	    Z                    ~� ��                          �� ��                         �� �C	    0                    �� ��                         �� ĕ                         � �D	    0                    0� ��                         N� Е                         l� `C	    P                    �� ��                         �� ܕ                   �            ��  C	    6                    �� ��                          � �                         $� �D	    P                    A� �                         _� ��                         }� @D	    6                    ��  �                          ��  �                         �� �#                          �� �#                          �  �                          G� 0�         w� ��         �� �         �� P�     .text   �                       .data                           .bss    P                            ��  �    N                   � (�                          V� �                         �� 0�    �                    �� @�                          �� �                         2� ��    ,                    [� T�                         �� $�                         �� �    $                    �� t�                         ڼ       0�                         2� P�    �                    `� ��                          �� <�                         �� p�                          �� С         � p�         G� Х     .text   �                       .data                           .bss    P                            v� p�    #                    �� ��                          �� H�                         � С                        F� ��                          |� T�                         �� p�    #                    �� ��                          � `�                         M� Х                        �� ��                          �� l�                         �� �                          � `�         :� ��         _�  �     .text   �                       .data                           .bss    P                            �� �    #                    �� ��   �                             �� x�                         	� `�                        6� ��                          d� ��                         �� ��    #                    �� ��                          �� ��                         �  �                        B� ��                          p� ��                         �� �X	                          �� pX	         �� ��                        
� ��         6�  �                        h�  �     .text   �                       .data                           .bss    P                            �� �X	    L                    �� ��                          �� ��                         �� pX	    D                    � ��                          B� ��                         j� ��                         �� ��                        �� ��                         � ̖                        �      6� �1                          I� �(         Y� `�	         �� `�         �� ��     .text   �                       .data                           .bss    P                             � �1    j                   � ��     l                    3� ؖ                         M� �(    t                   c� h�     T                    z� �                         �� `�	    '                   �� ��     p                    � �                         Y� `�    Y                   �� ,�     l                    �� ��                         � ��    Z                   L� ��     T                    �� �                         } �                         �� ��                          �� ��	         � 0�	     .text   �                       .data                           .bss    P                            ;� ��    �                     u� ��  �                              �� �                         �� ��	    �                     � ��                          B�  �                         n� 0�	                        �� ��                          �� ,�                     .rdata  �     �                     �� �                         	� �                         /�                           Q� @W                          � �!     p                    ��  !     p                    �� ��                          5� ��     .text   �                       .data                           .bss    P                            �� ��    /                    �� ��                          >� 8�                         �� ��    0                    �� �                          N� D�                         �� p                          �� �     .text   �                       .data           �                      .bss    P                            � p                        /� �                          X� P�                         �� �                        �� �                          � \�                         I� `�    *                   �� `�                          � ��    T                   �� ��         �� p�    !                   S� p�         �� @�    C                   .� @�         �� 0�    6                   � 0�         m�  �    V                   ��  �         M� ��    I                   �� ��         +� ��    q                   �� ��         �  �                       w�  �         �� `�    V                   U� `�         �� P�    V                   7� P�         �� ��    V                   � ��         �� p�    V                   � p�         }�  �    -        �                 ��  �         I� 0�    S                   �� 0�         � �    $                   �� �         �� ��    I                   b� ��         �� ��    9                   <� ��         �� @�    \                   � @�         �� ��    O                   �� ��         _�  �    w                   ��  �         ;  ��                       �  ��          ��    b                   � ��         � ��    b                   k ��         � �    b                   M �         � ��    b                   9 ��         �  �	     .text   �                       .data                           .bss    P                             �                         m h�                        � (�                         D t�                        � 4�                          ��                    �      .rdata  �     O                     � <�                          ��                        w D�                         � ��                        O	 P�                         �	 ��                        7
 X�                         �
 ��                         `�                         � ��                         p�                         r ȗ                        � t�                         X ԗ                        � |�                         B ��                        � ��                         , �                        � ��                           ��                        � ��                         	 �                        s ��                         � �                        M ��                         � �                        ' ��                         � �      (�                         ��                          4�                        � ��                         _ @�                        � ��                         F L�                        � ��                         + X�                        � ��                          d�                         ��                         � p�                        i ��                         � |�                        S ��                         � ��                        = �                         � ��                        ;  �	    *                    � �                         � ��                         E �                          ` @;         } Ф         � ��     (                   � Ф         � �         � ��     (                   � �          �C         . ��     �      (                   N �C         j ��         �  �     (                   � ��         � `�         � P�     (                   � `�          ��          ��         1 �C         M p�         e 0�         } ��         � ��     (                   � ��         � p�         � �         � ��     (                     �         .  ��         E  �         _  ��     (                   }  �         �  p         �  �7         �  0�     (                   �  �7         ! �7         !! p�         ;! p�         U! ��         p! ��         �! �C         �! �C         �! P�         �! P�         �! �         " �         5" 0�         Q" 0�         m" ��         �" ��         �" P         �" P         �" �7         �" �7     .text   �                       .data               �                  .bss    P                            # �                         8# ,�                          Z# ��                         |# @;                         �# 0�                          �# ��                         �# Ф    P                    $ 4�                          "$ Ę                         @$ �                        ^$ <�                          }$ И                         �$ �C                        �$ @�                          �$ ܘ                         % ��                        "% D�                          A% �                         `% `�                        ~% H�                          �% ��                         �% ��                        �% L�                          �%  �                         & ��    $                    3& T�                          R& �                 �              q& �C    $                    �& \�                          �& �                         �& p�    $                    �& d�                          ' $�                         5' 0�    $                    S' l�                          r' 0�                         �' ��    P                    �' t�                          �' <�                         �' p�                        ( |�                          /( H�                         O( �                        l( ��                          �( T�                         �( ��    $                    �( ��                          �( `�                         ) �                        !) ��                          B) l�                         c) p    $                    �) ��                          �) x�                         �) �7                        �      �) ��                          * ��                         ** �7    $                    K* ��                          m* ��                         �* p�    8                    �* ��                         �* ��                         �* ��                        + ��                          4+ ��                         V+ �C                        {+ ��                          �+ ��                         �+ P�                        �+ ��                          
, ��                         ,, �                        M, ��                          o, ̙                         �, 0�    8                    �, ��                         �, ؙ                         �, ��                        -  �                          :- �                         [- P                        ~- �                          �- �  �                             �- �7                        �- �                          . ��                         4. ��	                          �. ��	     .text   �                       .data                           .bss    P                            �. ��	                        0/ �                          �/ �                         �/ ��	                        :0 (�                          �0 �                         �0 �                          1 В         H1 �         r1 @�     .text   �                       .data                           .bss    P                            �1 �    �   
                 �1 8�     -                    2  �                     .rdata       �                    62 В    j  ,                 n2 h�                          �2 ,�                         �2 �    �   
                 3 p�     - �                         A3 8�                         r3 @�    j  ,                 �3 ��                          �3 D�                         4 P�                          64 pP                        Y4 P�         s4  �         �4 �         �4 Q                        �4 �         �4 ��         5 ��         5 ��         85 0�         R5 �P                        v5 0�         �5  C         �5 �Q                        �5  C         �5 �         6 �P                        26 �         L6 ��         f6 �P                        �6 ��         �6 p�         �6 p�         �6 @�         �6 �P                        7 @�         /7 �         K7 @Q                        q7 �         �7  7         �7 �Q                        �7  7         �7 ��         	8 ��         $8 p�         <8 p�         T8 `��               o8 `�         �8  �         �8  �         �8 P�         �8 P�         �8 �         9 ��         )9 ��         A9 �         [9 �         u9 е         �9 �P     .text   �                       .data                           .bss    P                            �9 P�                        �9 ��                         �9 P�                         :  �                        :: ��                         [: \�                         |: �                        �: ��                         �: h�                         �: ��                        ; ��                         ); t�                         L; ��    A                    k; ��                         �; ��                         �; 0�    !                    �; ��                          �; ��                         <  C    !                �          1< �                          V< ��                         {< �    !                    �< �                          �< ��                         �< ��    !                    �< �                          = ��                         ?= p�    A                    `= �                         �= ��                         �= @�    !                    �= 8�                          �= Ț                         > �    !                    %> @�                          H> Ԛ                         k>  7    !                    �> H�                          �> ��                         �> ��                        �> P�                          ? �                         ;? p�                        Y? T�                          x? ��                         �? `�                        �? \�                          �? �      �                         �?  �                        @ `�                          ?@ �                         a@ P�                        �@ h�                         �@ �                         �@ �                        �@ t�                         	A (�                         +A ��    4                    IA ��                          hA 4�                         �A �    %                    �A ��                         �A @�                         �A е                        	B ��                         *B L�                         KB �P    v                    zB ��                         �B X�                         �B ��                          C p�         3C `          hC P.          �C @�         �C @�          �C @�     __tcf_0  �	         D �         >D d	         `D  �     (             �            �D d	         �D �c	         �D p         �D �x         E p�     X   
                4E �x         SE �x         rE 0A         �E 0    2                   �E 0         �E ��     (                   F �    :                   6F �         OF ��         �F @�	         �F p^	         �F p^	         MG a	         �G a	         H  \	         OH  \	         �H ��	         �H �t                        �H ��                         �H �l                        I ��                         !I �t                        =I ��                         eI pq                        �I `c          �I ��          �I ��                         �I `�                         J �z     (               .text   �                       .data                           .bss    P                        .rdata  �     >                     @J�       ��                        sJ ��                          �J d�                         �J p�    T   	                 K ��                          @K p�                         sK @�                        �K ��                          �K |�                         �   �	                        �  ��                          	  ��                         L �    $                    1L ��                          aL ��                         �L d	                        �L ��                          �L ��                         M �c	    $                    3M ��                          \M ��                         �M p                        �M ��                          �M ��                         N �x                        0N ��                          VN ě                         |N �x    $                    �N ��   �                             �N Л                         �N 0A    E                    CO  �                          �O ܛ                         �O �                        P �                        1P �                        QP ��                        qP ��    �                    �P ,�                         �P  �                         *Q @�	                        IQ L�                          iQ �                         �Q p^	    �                   �Q T�     O                    DR �                         �R a	    �                   S ��     U                    }S $�                         �S  \	    o                   %T ��     >                    `T 0�                         �T ��	    h                   �T <�     I                    �T <�                         U `c                         5U ��     %   �                        dU @�     P   	                 �U `                          �U P.                         V  �                          SV  �         �V ��         �V ��         ;W `�         �W `�         �W PC         &X PC         wX  �         �X  �         Y �         ^Y �         �Y p�         �Y p�         CZ           �Z           �Z P7         1[ P7         �[ @�         �[ @�     .text   �                       .data                           .bss    P                            \  �    C                    m\ ��                         �\ H�                         ] ��    C                    g] ��                         �] T�                         ^ `�    !                    d^ ��                          �^ `�                         _ PC    !                    c_ ��                          �_ l�  �                             `  �    !                    f` ��                          �` x�                         a �    !                    aa ��                          �a ��                         	b p�    !                    [b ��                          �b ��                         c      !                    Vc ��                          �c ��                         d P7    !                    Xd ��                          �d ��                         e @�                        Ye ��                          �e ��                         f ж                          f ж         1f ��         ~f ��         �f `�         �f `�         g ��         g ��         7g ��         Rg �         jg �         �g �         �g �         �g �     .text   �                       .data                           .b�      ss    P                            �g ж                         �g ��                          h ��                         ,h ��                        h  �                          �h ̜                         'i `�                        Hi �                          ji ؜                         �i ��                        �i �                         �i �                         �i ��                        j �                         4j �                         Vj �                        tj $�                          �j ��                         �j �    K                     �j (�                          �j �                         k �    �                    4k ,�                         Uk �                         vk P�                          �k @�         �k �Q         l 0Q         Hl `�         ul `��               �l �         �l �     __tcf_0  �	         �l P�         +m и         Ym ��         qm ��     (                   �m ��         �m p�         �m @P         �m `�         )n `�     __tcf_1 0�	         dn PQ         �n П	         �n �          �n �z         o �z         )o �z         Go �z         do �          �o �z         �o ��         �o ��	         	p �c          6p `�          cp �c          �p  �          �p �          �p ��          q ��     P               .text   �                       .data                           .bss    P                        .rdata                             8q P�                        pq <�                          �q  �                         �q @�                        r @�                          Qr ,�                         �r �Q                         �r D�     �                           s 8�                         ?s 0Q                         ~s H�                          �s D�                         �s `�                         1t L�                          et P�                         �t �                         �t P�                          u \�                         �   �	                         �  T�                          	  h�                         7u P�                        ju X�                          �u t�                         �u и                        v \�                          ;v ��                         pv ��                        �v `�                          �v ��                         �v p�    $                    �v d�                          	w ��                         (w @P    e                    ^w l�                          �w ��           �                    �w `�    K                    x ��                          Qx ��                         �x 0�	                         �x ��                          �x ��                         �x PQ    [                    y ��                          Iy ȝ                         �y П	    �                    �y ��     !                    �y ԝ                         �y �z                         z ��                          ?z ��                         dz �z                        �z ��                          �z �                         �z �z                        �z ��                          { ��                         ={ �z                        a{ ��                          �{ �                         �{ ��    H                    �{ ��                          | �                         I| ��	                   �            �| ��                          �| �                     .ctors  `�	                        �| �c                         *} `�     *                     ^} �c                         �}  �     )                     �} �     P   	                 �} ��     P   	                 +~ �                         _~ �                         �~ P&                          �~ 0�     .text   �                       .data                           .bss    P                            �~ P&    z                   �~ ��     P                     (�                          0�    |                   P 8�     P                    � 4�                         } �                         � �I                          � �y         � ��     (                   ,� �y         L� �y     .text   �                       .data                           .bss  �        P                        .rdata  0                          l� �I                        �� ��                          �� @�                         � �y                        � ��                          9� L�                         `� �y    )                    �� ��                          �� X�                         ԁ �                           ��            �� p          	� �          � �          )� @	          <� �	          M� �	          ^� P
          l� �          w�           ��  ,          ��            �� �          �� �          ˂ `          � �          � �          � @          =�           L� �          [� @          f� �          x�       d_name  @      d_type  �           �� �6          �� ��	         �� �*          ă @/          ݃ �,          � p-          �� �/          �  0   �             � �0          0� �*          ;�  5          F� �;          Y� ~          f� �~          r� ��          �� ��          ��  �          �� ��          ̄ @�          ܄ P�          � ��          #� �          2� p�      .text   �     �  �             .data                           .bss    P                        .xdata  ��     @                .rdata  `     �  H            .pdata  d�       �                 P� ��	    �                     _� ��                          o� t�                         � `�	                      .text   ��                       .data                           .bss    P                            �� `�	    4                    �� ��                          ˅ ��                         � ��	                      .text   ��                       .data                           .bss    P                            � ��	    7   �                       '� ��                          K� ��                         o� P�	                      .text   ��                       .data                           .bss    P                            �� P�	    X                    �� �     $                    �� ��                         } �                         ӆ `                          � �d	         � 0�     (                   .� �d	         I� pd	         d�  d	         ��  d	         �� P�	         Ç ��	         �  �	         #� �q                        D� ��                     .text   ��                       .data                           .bss    P                            e� `                         �� (�                          �� ��                         ֈ �d	    P                    �� ,�                          � ��                         ;� pd	              �                \� 4�                          ~� ��                         ��  d	    H                    ĉ <�     %                    � Ƞ                         � P�	    V                    7� d�                          a� Ԡ                         �� ��	                         �� p�                          Ԋ �                         ��  �	                        A� t�                          �� �                     .file   _j  ��  ggccmain.c             Ӌ ��                       p.93846            � ��          �� �S                    __main  P�          � P       .text   ��     �                .data                         .bss    P                       .xdata  x�                      .pdata  ��     $   	             .file   gj  ��  gnatstart.c        .text   p�                       .data                           .bss    `                        .f�      ile   oj  ��  gwildcard.c        .text   p�                       .data   0                       .bss    `                        .file   j  ��  gcharmax.c              � p�                       .text   p�                     .data   @                       .bss    `                       .xdata  ��                      .pdata  �                     .CRT$XIC(                      .file   �j  ��  gdllargv.c         _setargv��                       .text   ��                      .data   P                        .bss    p                        .xdata  ��                      .pdata  (�                     .file   �j  ��  ggs_support.c          .� ��                           E� �.                         ]� �.                         �� p�          �� �           �� `          ��  ;      .text   ��     �               .data   P                        .bss    �      x                .xdata  ���                             .pdata  4�                     .rdata   ;                     .file   �j  ��  g_newmode.c        .text   p�                       .data   P                        .bss                           .file   �j  ��  gtlssup.c              ̌ p�                           ی ��          � �H                    __xd_a  `       __xd_z  h           �  �      .text   p�     �                .data   P                        .bss                          .xdata  ��                      .pdata  L�     $   	             .CRT$XLDH                      .CRT$XLC@                      .rdata   ;     H                .CRT$XDZh                       .CRT$XDA`                       .CRT$XLZX                       .CRT$XLA8                       .tls$ZZZ   	                    .tls        	                    .file   �j  ��  gcinitexe.c        .text   0�                       .data   P      �                        .bss                            .CRT$XCZ                       .CRT$XCA                        .CRT$XIZ0                       .CRT$XIA                       .file   �j  ��  gmerr.c                � 0�                           #�            1� ��      _matherr��      .text   0�     \               .data   P                        .bss                           .xdata  ��     $                 .pdata  p�     $   	             .rdata  �;     @               .file   k  ��  gCRT_fp10.c        _fpreset��                       fpreset ��      .text   ��                      .data   P                        .bss    0                       .xdata  ��                      .pdata  ��                     .file   k  ��  gmingw_helpers.c       H� ��                           X� ��      .text   ��                      .data   P                        .bss    0                      .xdata  �      ��                      .pdata  ��                     .file   3k  ��  gpseudo-reloc.c        h� ��	                          w� ��          �� D      the_secsH          �� ��          �� @           �S                        �  T                    .text   ��     �  $             .data   P                        .bss    @                      .rdata  �<                         P� ��	    i                    _�  �                          o� ��                     .xdata  �     (                 .pdata  ġ                     .file   ;k  ��  gxtxtmode.c        .text   P�                       .data   P                        .bss    P                      .file   Pk  ��  gcrt_handler.c          � P�                           :� �          P� h          _� �          i� �          s� �      .text   P�     w               .data   P                        .bss    `     �      �                .xdata  4�                       .pdata  ܡ     $   	             .rdata  �=                      .file   dk  ��  gtlsthrd.c             �� Ы                           ��  	          ��  	          Ǝ @�          � 	          �� ��          � `�      .text   Ы     j  '             .data   P                        .bss     	     H                 .xdata  T�     0                 .pdata   �     0                .file   lk  ��  gtlsmcrt.c         .text   @�                       .data   P                       .bss    `	                       .file   tk  ��  g    *�           .text   @�                       .data   `                        .bss    `	                      .file   �k  ��  gpesect.c              >� @�                           X� `�          k� ��          z� Ю          �� `�          �� �          ď  �          ׏ ��          � а          � p�      .text �        @�     �  	             .data   `                        .bss    p	                       .xdata  ��     H                 .pdata  0�     x                .file   �k  ��  gfake                  �  ��    .                    �                            �       {                .text    �     2                 .data   `                        .bss    p	                           �  `   
   0                    �       �                     �  H     H                .file   �k  ��  glibgcc2.c         .text   `�                       .data   `                        .bss    p	                           �  ��    �                   �       5                    �  �   
                        �  �     �                .file   �k  ��  gunwind-seh.c          &� `�                           B� ��          P� �          ^�  �          m� �          {�  �          �� 0�          �� @�   �             �� P�          Ґ `�          � ��          � ��          � ��          4� ��          K� �          Z� ��          t� �          �� �          �� 0�      .text   `�     '               .data   `                        .bss    p	                       .xdata  ��     �                 .pdata  ��     �   9                 �  ��    ;s  �                 �  O     ~                    ��        c                    �  �   
   0                    �  5     X                   �  �     �                     �  �     �  &             .file   l  ��  gemutls.c              �� ��                           ͑ и          ّ �	          � �	          � �          � p	          � x	          � �      .text   ��     z               .data   `                        .bss    p	                       .xdata  `�     (                 .pdata  ��     0                    �      �  �b    T(  �                 �  �     �                    �� c     N  	                 �  �   
   0                    5�        �                    �  �     �                   �  [     �                     �  x     �                .file   l  ��  gstrtodnrp.c       __strtod�                       fpi.4260`           C� �      .text   �     �                .data   `                       .bss    �	                       .xdata  ��                      .rdata  �=                     .pdata  ��                     .file   &l  ��  gstrtof.c          __strtof �                           R� �           \�  �      .text    �     �                .data   �                       .bss    �	                       .xdata  ��                      .rdata   >                     .pdata  ȣ                     .file   4l  ��  gbtowc.c           btowc   ��                       .text   ��  �         P                .data   �                        .bss    �	                       .xdata  ��                      .pdata  ԣ                     .file   Hl  ��  gmbrtowc.c             k�  �                       mbrtowc ��          x� �	          �� �          �� �	      mbrlen  �          �� �	      .text    �     8               .data   �                        .bss    �	                      .xdata  ��     @                 .pdata  �     0                .file   Pl  ��  gmingw_matherr.c   .text   @�                       .data   �                       .bss    �	                       .file   cl  ��  gstrtold.c             �� @�                       __eone  �>      __etens @>      strtold ��      .text   @�     �	  %             .data   �                        .bss    �	                       .rdata   >     �                 .xdata  ��     (                 .pdata  �                     .f�      ile   sl  ��  gwcrtomb.c             ˒ ��                       wcrtomb P�          ؒ ��      .text   ��     �               .data   �                        .bss    �	                       .xdata  �     (                 .pdata  (�     $   	             .file   �l  ��  gwctob.c           wctob   ��                       .text   ��     w                .data   �                        .bss    �	                       .xdata  0�                      .pdata  L�                     .file   �l  ��  gwctype.c          wctype  �                       cmap    `?      .text   �     `                .data   �                        .bss    �	                       .rdata   ?                    .xdata  8�                      .pdata  X�                     .file   �l  ��  gfopen64.c         fopen64 p�                       .text   p�                     .data   �                        .bss    �	               �              .xdata  D�                      .pdata  d�                     .file   �l  ��  gfseeko64.c        _flush  ��                       fseeko64�          � ��          � `T                        �  �          � ��          %�  @      .text   ��     �               .data   �                        .bss    �	                       .xdata  H�     H                 .pdata  p�     <                .rdata   @     p                .file   �l  ��  gftello64.c        ftello64`�                       .text   `�     )                .data   �                        .bss    �	                       .xdata  ��                      .pdata  ��                     .file   �l  ��  glseek64.c         lseek64 ��                       .text   ��                     .data   �                        .bss    �	                       .xdata  ��                      .pdata  ��                     .file   �l  ��  g�      mingw_vsnprintf.c     2� ��                       .text   ��     \                .data   �                        .bss    �	                       .xdata  ��                      .pdata  Ĥ                     .file   �l  ��  gstrtodg.c             D�  �                       rvOK    ��          T� @�          d� p�          s�  �          }� �T                        �� �B          �� T                        �� �T                    .text    �     J   l             .data   �                        .bss    �	                       .xdata  ��     T                 .pdata  Ф     <                .rdata  �A     �  .             .file   
m  ��  gsum.c                 ܓ P�                       .text   P�     H               .data   �                        .bss    �	                       .xdata  ��                      .pdata  �                     .file   %m  ��  gcephes_emath.c    __m16m  �      ��                           � P�      __emovi @�      __eaddm  �      __esubm `�      __edivm ��      __emulm  �      __toe64 @�      __ecmp  ��      __eshift��          �� ��           � ��      __emovo �     __emul  P     .text   ��     [                .data   �                        .bss    �	                       .xdata  �     �                 .pdata  �     �   *             .file   Em  ��  gmingw_pformat.c       
�                        fpi.6121�           � �         '� P         ;� `	         N� 0
         ]� �
         w�           ��           �� �         �� �         ̔ p         � P         �           � �         �           -�       .text        !  !             .data   �                       .bss    �	                       .xdata  ��     �                 .pdata  ��     �   0             .rdata   C     �  [           �        .file   Vm  ��  gdmisc.c               =� (                          L� @(         \� �(         g� �(     .text   (    |               .data   �                        .bss    �	                       .xdata  ��     0                 .pdata  ��     0                .file   fm  ��  ggdtoa.c           __gdtoa �*                      .text   �*    �  Q             .data   �                        .bss    �	                       .rdata  �D     �                .xdata  ��                      .pdata  ��                     .file   vm  ��  ggethex.c              t�  @                          �� 0T                    .text    @    	               .data   �                        .bss    �	                       .xdata  ��                      .pdata  ��                     .file   �m  ��  ggmisc.c               �� 0I                          �� 0J     .text   0I    C                .data �        �                        .bss    �	                       .xdata  ��                      .pdata  Ȧ                     .file   �m  ��  ghd_init.c             �� �J                      .text   �J    �                .data   �                        .bss    �	                       .rdata  PE                      .xdata  �                      .pdata  �                     .file   �m  ��  ghexnan.c              ϕ  K                      .text    K    �               .data   �                        .bss    �	                       .xdata  �                      .pdata  �                     .file   �m  ��  gmisc.c                ܕ �N                          �           �             � �O         � �O     freelist�          � �           )� �	          5� �P         A� PQ         O�  R         Y� 0R         d� `S     p5s     �	          s� �E          }� �T  �             �� �U         ��  V         �� �W         �� �X         �� �Y     .text   �N    #  +             .data   �                      .bss    �	     �	                .xdata  (�     �                 .pdata  ��     �   *             .rdata  �E     H                .file   �m  ��  gsmisc.c               �� �Y                          ɖ �Z         Ֆ �[         � �[         � @\     .text   �Y    �               .data   �                        .bss    �                       .xdata  ��     4                 .pdata  ��     <                .file   �m  ��  gstrnlen.c         strnlen �\                      .text   �\    (                 .data   �                        .bss    �                       .xdata   �                      .pdata  ܧ                     .file   �o  ��  gwcsnlen.c         wcsnlen ]                      .text   ]    !                 .data   �          �                    .bss    �                       .xdata  �                      .pdata  �                     .text   @]     .data   �       .bss    �      .idata$7�      .idata$5	      .idata$4�      .idata$6:      .text   H]     .data   �       .bss    �      .idata$7|      .idata$5	      .idata$4�      .idata$60      .text   P]     .data   �       .bss    �      .idata$7x      .idata$5�      .idata$4�      .idata$6$      .text   X]     .data   �       .bss    �      .idata$7t      .idata$5�      .idata$4�      .idata$6      .text   `]     .data   �       .bss    �      .idata$7p      .idata$5�      .idata$4|      .idata$6      .text   h]     .data   �       .bss    �      .idata$7l      .idata$5�      .idata$4t      .idata$6      .text   p]     .data   �       .bss    �      .idata$7h      .idata$5�      .idata$4l      .idata$6�      .text   x] �          .data   �       .bss    �      .idata$7d      .idata$5�      .idata$4d      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7`      .idata$5�      .idata$4\      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7\      .idata$5�      .idata$4T      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7X      .idata$5�      .idata$4L      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7T      .idata$5�      .idata$4D      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7P      .idata$5�      .idata$4<      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7L      .idata$5�      .idata$44      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7H      .idata$5�      .idata$4,      .idata$6�      .text   �]     .d�      ata   �       .bss    �      .idata$7D      .idata$5�      .idata$4$      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7@      .idata$5�      .idata$4      .idata$6�      .text   �]     .data   �       .bss    �      .idata$7<      .idata$5�      .idata$4      .idata$6�      .text   �]     .data   �       .bss    �      .idata$78      .idata$5|      .idata$4      .idata$6z      .text   �]     .data   �       .bss    �      .idata$74      .idata$5t      .idata$4      .idata$6p      .text   �]     .data   �       .bss    �      .idata$70      .idata$5l      .idata$4�      .idata$6d      .text   �]     .data   �       .bss    �      .idata$7,      .idata$5d      .idata$4�      .idata$6Z      .text   �]     .data   �       .bss    �      .idata$7(      .idata$5\      .idata$4�      .idata$6R      .text   �]     .data   � �            .bss    �      .idata$7$      .idata$5T      .idata$4�      .idata$6J      .text    ^     .data   �       .bss    �      .idata$7      .idata$5D      .idata$4�      .idata$66      .text   ^     .data   �       .bss    �      .idata$7      .idata$5<      .idata$4�      .idata$6,      .text   ^     .data   �       .bss    �      .idata$7      .idata$54      .idata$4�      .idata$6"      .text   ^     .data   �       .bss    �      .idata$7      .idata$5,      .idata$4�      .idata$6      .text    ^     .data   �       .bss    �      .idata$7      .idata$5$      .idata$4�      .idata$6      .text   (^     .data   �       .bss    �      .idata$7      .idata$5      .idata$4�      .idata$6      .text   0^     .data   �       .bss    �      .idata$7       .idata$5      .idata$4�      .idata$6�      .text   8^     .data   �       �      .bss    �      .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   @^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4�      .idata$6�      .text   H^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4�      .idata$6�      .text   P^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4|      .idata$6�      .text   X^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4t      .idata$6�      .text   `^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4l      .idata$6�      .text   h^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4d      .idata$6�      .text   p^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4\      .idata$6�      .text   x^     .data   �       .bss    �      �      .idata$7�      .idata$5�      .idata$4T      .idata$6�      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4L      .idata$6�      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4D      .idata$6�      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4<      .idata$6~      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$44      .idata$6v      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4,      .idata$6l      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4$      .idata$6b      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5�      .idata$4      .idata$6X      .text   �^     .data   �       .bss    �     �       .idata$7�      .idata$5�      .idata$4      .idata$6P      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5|      .idata$4      .idata$6F      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5t      .idata$4      .idata$6>      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5l      .idata$4�      .idata$64      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5d      .idata$4�      .idata$6*      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5T      .idata$4�      .idata$6      .text   �^     .data   �       .bss    �      .idata$7�      .idata$5<      .idata$4�      .idata$6�      .text   �^     .data   �       .bss    �      .idata$7�      .idata$54      .idata$4�      .idata$6�      .text   �^     .data   �       .bss    �      .idata�      $7�      .idata$5,      .idata$4�      .idata$6�      .text    _     .data   �       .bss    �      .idata$7�      .idata$5$      .idata$4�      .idata$6�      .text   _     .data   �       .bss    �      .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   _     .data   �       .bss    �      .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   _     .data   �       .bss    �      .idata$7|      .idata$5      .idata$4�      .idata$6�      .text    _     .data   �       .bss    �      .idata$7x      .idata$5�      .idata$4�      .idata$6�      .text   (_     .data   �       .bss    �      .idata$7t      .idata$5�      .idata$4�      .idata$6�      .text   0_     .data   �       .bss    �      .idata$7p      .idata$5�      .idata$4|      .idata$6�      .text   8_     .data   �       .bss    �      .idata$7h   �         .idata$5�      .idata$4l      .idata$6l      .text   @_     .data   �       .bss    �      .idata$7`      .idata$5�      .idata$4\      .idata$6L      .text   H_     .data   �       .bss    �      .idata$7X      .idata$5�      .idata$4L      .idata$6.      .text   P_     .data   �       .bss    �      .idata$7T      .idata$5�      .idata$4D      .idata$6      .text   X_     .data   �       .bss    �      .idata$7P      .idata$5�      .idata$4<      .idata$6      .text   X_     .data   �       .bss    �      .idata$7L      .idata$5�      .idata$44      .idata$6       .text   `_     .data   �       .bss    �      .idata$7D      .idata$5�      .idata$4$      .idata$6�      .text   `_     .data   �       .bss    �      .idata$7@      .idata$5�      .idata$4      .idata$6�      .text   h_     .data   �       .bss    �      .idata$7<      .ida�      ta$5�      .idata$4      .idata$6�      .text   p_     .data   �       .bss    �      .idata$78      .idata$5|      .idata$4      .idata$6�      .text   x_     .data   �       .bss    �      .idata$74      .idata$5t      .idata$4      .idata$6�      .file   	p  ��  gacrt_iob_func.c       �� �_                      .text   �_                    .data   �                      .bss    �                       .xdata  �                      .pdata  ��                     .file   p  ��  g    ��               � �_                      handler �          1� �_         P� �_         t� �_     .text   �_                    .data   �                      .bss    �                      .xdata  �                      .pdata   �                     .file   +p  ��  g__p__acmdln.c         �� �_                          �� pT                    .text   �_              �            .data                         .bss    �                       .xdata  �                      .pdata  �                     .file   ;p  ��  g__p__fmode.c          ؗ �_                          � �T                    .text   �_                    .data                        .bss    �                       .xdata  �                      .pdata  $�                     .file   Wp  ��  gfake              hname         fthunk  t      .text   �_                      .data                           .bss    �                       .idata$2                      .idata$4      .idata$5t      .text   �_     .data          .bss    �      .idata$7\      .idata$5�      .idata$4T      .idata$6B      .text   �_     .data          .bss    �      .idata$7H      .idata$5�      .idata$4,      .idata$6�      .file   ep  ��  gfake              .text   �_                      .d�      ata                           .bss    �                       .idata$4�                      .idata$5	                      .idata$7�                      .file   �p  ��  gcond.c                �� �_                          � �`     fo      �           � �          ,� �`         7� pa         P� �a         f� �a         �� �a         �� �a         �� b         И �b         � �b         �� d         �            � pd         1� @g         @� �g         U� pi         i� �j         �� �k         �� @m         �� �n         �� pp         ҙ �p     .text   �_    �  Z             .data                          .bss    �                      .xdata   �     �                 .pdata  0�       B             .rdata  �F     "                 .file   �p  ��  gmisc.c                �� �p                          	� �p         +� q     .text   �p�          �                .data   0                       .bss    �                       .xdata  �                      .pdata  8�     $   	             .file   �p  ��  gmutex.c               C� �q                          S�  r         f� 0s         ~� �t         �� `u         �� �u         �� 0v         Қ pv         � �v         � �v         � �v         7� �v         T�  w         q� 0w         �� @w         �� `w         Λ pw     .text   �q    �               .data   0                       .bss    �                       .xdata  0�     x                 .pdata  \�     �   3             .file   �p  ��  gspinlock.c            � �w                          � �w         � �w         (� �w         =� �w     .text   �w    j                 .data   0                       .bss    �                       .xdata  ��                      .pdata  (�     �      <                .file   7q  ��  gthread.c              Q� �w                          c� x         s� 0      once_obj�          � �x         �� H          �� �x         �� �      idList  �          �� `y         ؜ �          � �          � �z         � 8          � �          !� �          +� @|         B�  }         X� 0}         h� �}         �� �~         ��            �� @         ӝ ��         � Ѐ         � @          � ��         *� �          C� ��         Z� ��     .tl_end (�         d� ��          � �          u� Ѕ         �� ��         �� ��         �� ��         ؞ `�         � ��         �� �          	� �          �  �         -�  �         A� p�         U� p�         c� ��         y� ��         �� ��         �� ��         ��  �         �� @�         ҟ           � �      P�         �� `�         � `�         �           1� ��         E� Ў         \� 0�         o� ��         ��  �         �� ��         �� 0�         ��  �         à ��         ֠ ��         � Г         ��  �         � 0�         ,� P�         H� `�         e� ��         �� ��         �� ��         �� Д         ȡ ��         � �         ��  �         � �         -� ��         C� �         R� ��         _� ��         p� �         � �         �� �          ��  �         Ţ 0�         آ 0�     .text   �w    E&  D            .data   0                      .bss    �     l                 .xdata  ��     �               .pdata  d�     0  �             .rdata  G     �                 .CRT$XLFP                      .file   �r  ��  grwlock.c              � @�                          �� X          � ��    �           � @�         ,� ��         C� ��         R�  �         \� ��          �           j� ��         t� @�         ��  �         � P          �� ��         �� �         �� У         ף p�         �  �         � ��         $� p�         :� �         P�  �         k� ��         �� ��         �� �         ��  �     .text   @�    �  Z             .data   P                      .bss                          .xdata  l�                     .pdata  ��       E             .rdata  �G     �                 .text    �     .data   `      .bss           .idata$7      .idata$5\      .idata$4�      .idata$6n      .text   (�     .data   `      .bss           .idata$7      .idata$5T      .idata$4�      .idata$6X      .text   0�     .data   `      .bss           .idata$7      .idata$5L      .idata$4�      .idata$6>      .text �        8�     .data   `      .bss           .idata$7      .idata$5D      .idata$4�      .idata$6.      .text   @�     .data   `      .bss           .idata$7      .idata$5<      .idata$4�      .idata$6      .text   H�     .data   `      .bss           .idata$7      .idata$54      .idata$4�      .idata$6       .text   P�     .data   `      .bss           .idata$7      .idata$5,      .idata$4�      .idata$6�      .text   X�     .data   `      .bss           .idata$7       .idata$5$      .idata$4�      .idata$6�      .text   `�     .data   `      .bss           .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   h�     .data   `      .bss           .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   p�     .data   `      .bss           .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   x�  �         .data   `      .bss           .idata$7�      .idata$5      .idata$4�      .idata$6�      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4|      .idata$6`      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4t      .idata$6L      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4l      .idata$62      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4d      .idata$6"      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4\      .idata$6      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4T      .idata$6      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4L      .idata$6�      .text   ��     .dat�      a   `      .bss           .idata$7�      .idata$5�      .idata$4D      .idata$6�      .text   ��     .data   `      .bss           .idata$7�      .idata$5�      .idata$4<      .idata$6�      .text   Ȫ     .data   `      .bss           .idata$7�      .idata$5�      .idata$44      .idata$6�      .text   Ъ     .data   `      .bss           .idata$7�      .idata$5�      .idata$4,      .idata$6�      .text   ت     .data   `      .bss           .idata$7�      .idata$5�      .idata$4$      .idata$6�      .text   �     .data   `      .bss           .idata$7�      .idata$5�      .idata$4      .idata$6p      .text   �     .data   `      .bss           .idata$7�      .idata$5�      .idata$4      .idata$6\      .text   �     .data   `      .bss           .idata$7�      .idata$5|      .idata$4      .idata$6J      .text   ��     .data   `  �          .bss           .idata$7�      .idata$5t      .idata$4      .idata$60      .text    �     .data   `      .bss           .idata$7�      .idata$5l      .idata$4�       .idata$6      .text   �     .data   `      .bss           .idata$7�      .idata$5d      .idata$4�       .idata$6      .text   �     .data   `      .bss           .idata$7�      .idata$5\      .idata$4�       .idata$6�
      .text   �     .data   `      .bss           .idata$7�      .idata$5T      .idata$4�       .idata$6�
      .text    �     .data   `      .bss           .idata$7�      .idata$5L      .idata$4�       .idata$6�
      .text   (�     .data   `      .bss           .idata$7�      .idata$5D      .idata$4�       .idata$6�
      .text   0�     .data   `      .bss           .idata$7�      .idata$5<      .idata$4�       .idata$6�
      .text   8�     .data   `      .b�      ss           .idata$7�      .idata$54      .idata$4�       .idata$6�
      .text   @�     .data   `      .bss           .idata$7�      .idata$5,      .idata$4�       .idata$6p
      .text   H�     .data   `      .bss           .idata$7�      .idata$5$      .idata$4�       .idata$6V
      .text   P�     .data   `      .bss           .idata$7x      .idata$5      .idata$4�       .idata$6*
      .text   X�     .data   `      .bss           .idata$7t      .idata$5      .idata$4�       .idata$6
      .text   `�     .data   `      .bss           .idata$7p      .idata$5      .idata$4�       .idata$6
      .text   h�     .data   `      .bss           .idata$7l      .idata$5�      .idata$4�       .idata$6�	      .text   p�     .data   `      .bss           .idata$7h      .idata$5�      .idata$4�       .idata$6�	      .text   x�     .data   `      .bss                  .idata$7d      .idata$5�      .idata$4|       .idata$6�	      .text   ��     .data   `      .bss           .idata$7`      .idata$5�      .idata$4t       .idata$6�	      .text   ��     .data   `      .bss           .idata$7\      .idata$5�      .idata$4l       .idata$6�	      .text   ��     .data   `      .bss           .idata$7X      .idata$5�      .idata$4d       .idata$6�	      .text   ��     .data   `      .bss           .idata$7T      .idata$5�      .idata$4\       .idata$6l	      .text   ��     .data   `      .bss           .idata$7P      .idata$5�      .idata$4T       .idata$6X	      .text   ��     .data   `      .bss           .idata$7L      .idata$5�      .idata$4L       .idata$6H	      .text   ��     .data   `      .bss           .idata$7H      .idata$5�      .idata$4D       .idata$6:	      .text   ��     .data   `      .bss                 .idata$7D      .idata$5�      .idata$4<       .idata$6	      .file   s  ��  gmingw_getsp.S         ڤ ��                      longjmp ƫ     .text   ��                    .data   `                       .bss                            .text   Ы     .data   `      .bss           .idata$7       .idata$5L      .idata$4�      .idata$6@      .text   ث     .data   `      .bss           .idata$7      .idata$5      .idata$4�      .idata$6�      .text   ث     .data   `      .bss           .idata$7�      .idata$5\      .idata$4�      .idata$6       .text   �     .data   `      .bss           .idata$7�      .idata$5L      .idata$4�      .idata$6
      .text   �     .data   `      .bss           .idata$7�      .idata$5D      .idata$4�      .idata$6       .text   �     .data   `      .bss           .idata$7�      .idata$5      .idata$4�      .idata$6      �      .text   �     .data   `      .bss           .idata$7l      .idata$5�      .idata$4t      .idata$6v      .text   ��     .data   `      .bss           .idata$7d      .idata$5�      .idata$4d      .idata$6Z      .file   !s  ��  gcygming-crtend.c      � �	                      .text    �                      .data   `                       .bss                                �� �	                        � p�                          � ��                         &� h�	                        3� ��          W� `�          �� �           �� �          � �O          3�  u      setvbuf �]         ^� �Q          ~� ��          �� ��          ¦            ߦ @J          � �          � 0       fdopen  (_         '� ��          :� �b          ^� �l          �� �          �� Pz          �� �          ˧  �      memcmp  ^         ��  �                � @]          .� 0T      towupperx]         C�  T          i� ,          v� �P      _ZTVSo  0�          ��  u          ��  �          �� �V          ֨ ��          � pp          4� �          B� P�          ]�  ~          q� ��     abort   �^         }� �P          �� <          �� ��          �  �          � 0�          Q� ��          c� �H          �� z          �� ��          ͪ ��         ߪ �          � ��         	� x�         � �          *� �W      realloc �]         P�           ]� �          q� 8       write   �^         �� �          �� �          ū �{          � �          �             � y          7� D          J�           W� p�          �� @b          �� @U          Ѭ  W          � �I          � @L          .� �Y          O� W          h�  #          �� pN          �� �z          ��       `O          ۭ �E          � L          � @�         �  N          f�           �� `Y          �� �          �� ��          ʮ  �          ޮ �          � �^         �� �L          P� 	          \� PU          m� �y          �� 0\          �� ��         Ư �          ԯ P$          �� @d          *� ��          N� �          \� ��          q� p$          �� ��          �� `�          �� 0      _ZTVSd  `�          װ �          � �J          ;� �H          K� �m          o�            �� @#          �� �}          � ��          0�  �          L� �N          _� �#          �� x�         �� ��         ɲ c          � ��          �            c� �K          ��  �          �� @\          г �t          �           �� p          <� �$          R�  ^          l� �q          �� �          �� �      fgetpos �^               �� �R          ô �#          ش �u          � ��          B� �         a� �          �� �s          �� ��          Ե ��          � @          � `N          $� �I          K� pm          o� �          �� ��         ��             �� �          �� �}          Ҷ �$          � �          "� �w          =� L          J� @Q          i� �_          �� `L          �� PT          � ��          4� ��          Z� @M          �� �S          �� `�          ˸ ��      signal  �]         ۸ 0�          �� �Q          "� `�          <� �Y          \� ��          �� ��          �� ��          �� �          �� �      strcmp  �]         й @          ݹ  �          � P]          .� pM          X� 0�          �� �          �� �Q          ͺ �I          � ��          � �          $� l          =�    ��       R� �\                g� �          �� ��          �� �S          � �v          �  �          � �           D� pn          i�  �          �� `}          �� @T          ϼ `�          �� ��           �  M          i� `t          ~� `�          �� 4          ��  �      memset   ^         �  �          	� ��          4� �          U� �          a�  �          �� ��          ˾ �d          �� h_         �  �          �  �          ;�  �          Q� |          ^�           l� �N          ~� �Q          �� ��          ˿ ,          � �          � �M          L�     ��       ]� `U          n�    ��       �� @�          �� �W      Sleep   �          �� �"          	� �#          !� �          6�  ]          L� �U          f� ��          �� �J          �� @W      _fmode  P          �� ��          �� �      malloc  (^     __xc_a              � �S                S� <          f� �          u�  t          �� �z          ��  �          �� �          �� p]          �� �      SetEvent��         �  O          3� 4      wcscoll X]         @�  �          �� T          �� �]          �� 0          �� ��          �� ��          � @{          0� ت         ;� �a          �� 0P          �� �S          �� ��          � �          #�  �          D�             ]� `�      memmove ^         �� Ѐ          �� �"          �� �         �� �          � ��          *� `K          E�  I          q� p          �� ��          ��     ��       �� ��          �� �#          � Ps          1� �Q          V� p�         g� J      fflush  �^         �� @u      strncmp �]     wcsftimeP]         �� 0"          �� �.          �� p�          �� �K          � �          6�  [          J� �l                g� �          ~� �           �� �R          �� �Z          �� �K          �           #� �         4� �O          �� 0Q          �� `�          �� �J          �� �T           � �          -� ��          I�  �         Z� p�         k� �u          �� �$          ��           �� ��          �� �b          � \          9� P          |�           �� �V          �� �          �� `�     _ZTISo   r          �� @_         �� P�          �� `d          (� 0�          E� �V      _ZTISd  �q          ^� �          �� 0      strxfrm �]         �� X          �� `~          �� �[      _ZTISi  �q          �� $           � P_         &� �\          :� ��          g� �t          }� �I          �� n          �� `          � ,          � �P          8�  c          a�  �          �� P�          �� �r          �� �          �  	                � �R          4�  �         H� �          e� �          {� �[          �� �N      putwc   �]         �� Ц      fclose  �^         �� $          �� ��          �� ��          � @�          � �          &�  �          d� 0$          �� �M          �� �\          �� �          �� �"      _ZTSSi  Д          � `�          2� �d          _� ��          �� @I          �� �O      _ZTSSd  ��          �� ��          �� `P          � �$          N� �          s� `F      strdup  �         �� �T          ��  �          �� ��          ��  �          ��  �          � ��         6� �          a�            �� t          �� ��          �� �          �  !          A� �O          f� @�          ��           �� T          ��  J          �� ��          �� ��          #�  �          c� @&          m� �H          �� P#      
      _ultoa  ث         �� 	          �� ��          � 0          ;�  �      _ZTSSo  ��          W� 0�          �� �U          �� q          �� ��          �            $�  �          H� �T          [� �      vfprintf`]         y� @�      strcoll �]         ��  �          �� �m          �� `          �� �P          � `I          4� �#          K� @;          U� @_          �� P          �� 0�          �� T          �� �v           �  {          !� �          1� �          M� @N          �� 0          ��  �      __xc_z             ��  Z          ��  �          � �          (� @�          T� @S          �� ��          ��    	        �� ��         ��  K          �   @ ��       $� p#          o� 0�          �� 0K          �� `           �� p�          � �          #� (�         7� ��          M� `�          r�  �          ��        �         ��  O          �  �          L� �          e� �T          t� �          �� p"          ��           �� `�          ��           �� �          �� �)          �� ��          � ��          (� 0�          o� �M          �� PR          ��           � @          *� pw          A� pK          c� �          v� ��          �� T          �� �K      __xl_z  X           �� ��          �           "� �          :� �          `� У          s�  �          �� @Y          �� �K          �� ��         �� �V          �� �          � d          � �^          =� ��          �� `S          ��  L          �� �L      __xl_c  @           � pQ          `� t      __xl_d  H           l�  �          �� ��          �� ��          �� pV          �� ��          � �          � pL          l� @R          �� �          �� @~                �� \          �� �          �� �          	� �n          Z� x�	         i� �M          �� �x          ��  M      __xl_a  8           � ��          3� PL          Y� �"          v� �(      _onexit �^         �� 8      __xl_f  P           ��            �� ��          �� `�          � o          0� px          w� �~          ��            �� ^          �� �]          �� 0U          	� `�          4� Pn          Y�  Q          �� 	      printf  Ы         �� ��          �� ��          ��  �          �� p^          �� 8�         � �          ,� �          8� p\          L� ��          x� ��          �� ��          �� �~          +� `�          V� Pq          �� 0�          �� �t          ��            �� Ъ         �� �_         � ��          �  �      fwrite  `^         6� `          P� �          `� `          ��       �[          �� �           � ��          �  �          ?� �          J� Pr          ]� |          r� �w          �� l          �� ��         �� S          �� 0]          �� P�          � ��          a� ��          �� Q          �� @�          � �         � �          6� @}          [� L      getwc   H^         x� �I          �� p_         �� ��          �� �o          �� PN          .� @c          X� p�          �� ��          �� �M          �� �y          � �l          !� po          =� �.          Z� `�          n� `�          �� ��          �� 0m          �� �          �� PV          �� ,          � �          C� ��      _CRT_MT P       wcsxfrm @]         �� ��          �� \          �� ��          �� �$          �  }      fsetpos h^         1�  %          t� �          �� pr      TlsAlloch�         ��    ��             �� `�          ��  Z          ��            �    ��       -� 0q          w� �R          �� �S          �� p          �� ��          � ��          �  a          G� ��         ^�           ��  U          �� �          �� �o          �� �_          � �          ,� �          :�  ^          E�            U� ��          f�  �          �� U          �� X�         �� �          �� �p      exit    �^         �� ��          � �R          V�           n�             �� @          �� ��      fprintf �^         �� Py          �� `M          �� @|          � `Z          2� t          @� `          Y� �|          ~� (�         �� L          ��  �          �� ��          �  �          F� �N          [� ��          r� @�          ��     	        �� 0y          �� p�          �� �r          �� �s          �� ��                �  �          i� �c          �� �"          �� `�          �� �W          #� �          =� 0x          �� �I          �� PY          �� pJ          �� ��          ��     ��       � �          3� PJ          X� �n          }�  �          �� `_         �� pT          �� 0�          �� T          ��  �          �  �          d�             |� ��         �� �W          �� �x          �� �          �� ��          � `�          Q� ��          �� ��          �� Pp          	� �          �           -� �b          r� �          �� `�          �� �      __end__    	        �� `"          �� t          �� 0I          � �\          "� �          0� �p          z� x_         ��            �� �P          � ��          1� �          D�            V� �          a� �[          �� ��          �� �Z      strtoul �]         ��  ~                �� pU            ��          =   J          b  py          �  �L      fread   x^         �  pv           Pa          G `'          Q ��          v ��         � ��         � �I          � `T          � @�            $          0 �          P �$          � `�          �    ��       � pq          � �          � `{           ��          H @�          c p�          � ��          � �N          � |      wcslen  H]          `J          / �o          K �          X �x          t 0`          �  �          � @V            N          V  d          � d          � �O          � �N           pI          5 �          M  �          s d          � Px          � �            �      getchar P^         \ �]         f ��          � �L      calloc  �^         �  �          � D                 X_           _          ��          : �K          X            j @"      _write  �^         � ]          � ��          � @�          �  $          +	 �|          P	 �          r	  �          �	 �^         �	  U          �	 �          �	 0o          �	 �]          
 \          
 ��          4
 ��          Z
 @P          |
 4          �
    ��       �
 �w          �
 �F          �
 `�          �
 �            �          1 �K          V ��          { @t          �  �          � ��          �  �          � PM          " PK          = �          I  S          d �$          � `�          � `�          B 0�          S M          p �      read    �^         � v          �            � �          � �          � �y          � �J           `$          3  d          m �         � `                 � ��          � ��          �  "          � P�         � P          	 �                     (  R          R `           d ��          �  P          � `#          � 0w          �  �           `R      ungetwc h]         A �          T �T          u  P          � �          �  v      fputc   �^         � ��          � �          
 @�      _fstat64_         ) @�          h  V          � �          �     ��       �    ��       � Ȫ         � 0O           �          = �n          �  I          � �N          � P�      iswctype8^         � 0z           \           $          ;  �          y  �          � P�         � �}          � ��           �w          5 p�          t @          � �T          � �V          � `�         � 0J           ��          $ t                9 8           K �#          b x�	         p �          � �J          � �+          � �V           �           $          [ 0�         h �          � ��          � �O      _ZSt3cin %          � @�                     9             G @�         V P�          �           � �R          � �z          � �            \          ; ��          ]  T          } 0L          � ��          � �l          �     ��       � ��           PQ          D ��          h `Q          � �Q      towlower�]         � `           � �          �           �             �          F H�         _ @�          � �]          �           � p[          �  �          � `           � P"      fputs   �^          <          ( 0[          F �`          � ��          �  �          � 0          �           	                   Q @K          y @�          � ��          � ��           Pv          K �~          �  �          � �U          � �R           R          D �J          f �]          � ��          � ��          � @�          � �          	  �          P �Q          � N          � s          � ��          �  �          :  �\      _fileno _         N  $          `  �!          �  �~          �  (           �  �           �  �          ! �S          >!           I! (      _charmax@           c! �          n!  �          �! `W          �! pW          �!  �          �! �"          " �V          '"  �          H" �M          f" �          �" pS          �" <          �" �\          �" �T          �" �{          �" �          # p�          # �          (# ��          h# pz          �#                  �#  �	         �# H_         �# @�          �# �[          �# X�         $ �          $             +$ �[          Y$  X          z$  ]          �$ �]          �$ �"          �$ �P          �$  _         �$ �      _cexit  8_         % ��          L% ��          �% �          �% ��          �%  L          "& ��          ?& �          N& �a          �& ��      free    p^     strftime�]         �&  �          �& �          �& `          �& �.          �& 0�         ' ��          .' �          N' ��          {' ��          �' ��          �' �Q          �'  �	         �' �L          �' �          ( @          R( PI          (  Q          �( �          �( �          �( @�          )) `�          E) �\          Y) `u      _setjmp �         �)  $          �) �w          �) @�          
*           !*     ��       6*       �W          \*           s* 0n          �* I          �* l      ungetc  p]         �* �      _ZTTSi   �          �*  �          �*  K      _errno  0_         +  }          6+ w          R+ �L      memchr   ^         �+ �u          �+ �          �+ �s          ,  �          /, �$          r, �R          �,  X          �, �n          �, �#          -  �          V- �O      _ZTTSd  �          �-           �- ��          �- ��          . ��          $.  S          <. pP          X. ��          �. �L          �. �L      __dll__     ��       �. P[          /  -          / 0W          0/ ��          G/ pO          k/ ��          �/ 0p          �/ �\          �/ �          �/ �v          &0 ��          G0 ��          s0 PP          �0  �          �0 d          �0 �P          �0 ��          1 �U      strerror�]     fopen   �^               ,1 ��         >1 `�          n1 ��      isspace @^         �1 @O          �1 h�         �1 ��          �1  {          2 ��           2 ��          <2 �          W2 `�          �2 @      _ZTTSo  0�          �2 PS          �2 pR          �2 �[          3 ��          53 PW      _tls_end   	    fileno  _         T3 �#          i3 @[          3 �          �3 �          �3 �          �3 @$          �3 ��         4 0V          ?4 %          �4 0#          �4 �          �4 �J          �4 �         �4 @�      putc    �]         5 x          65   @ ��   sprintf �]         B5 �J          a5 0R          �5 0S      __xi_z  0           �5 �]          �5 �S          6 0�          M6    ��       `6 P\          s6 O          �6 �c      getc    X^         �6 ��          7 �N          D7 ��          j7 #      memcpy  ^               �7 �r          �7 �          �7 �"          �7 `V          �7 �t          8 �I          (8  R          R8 0N          �8 �          �8 �S          (9 0�          @9 ��          �9 ��          �9 �*          �9 �          �9 0v          �9 �P          : p�          /: �O          �: �M      strlen  �]         �:  �          �: @�          �: 0          B; �[          i; ��          �; PO          �; `\          �; ��          �; ��          �; $          < P          )< @�          C< |          P<  ;          h< `�          �< 0M          �< L          �< H�         �< 4          = �M          7=  �          X= �]          p=    ��       �=  #          �= ��         �= �s          �=            �=     ��       > �V          > �T          8> D          F> ��          {> �y          �> D          �>  �          �> �                �> `[          �> ��          ?  W          ? Po          G?  �      _ZTVSi  ��          l?  |          �?  \          �? �          �? `]          �? @�          �? ��          #@ `�          >@ K          b@ �x          z@ ��          �@ ��          �@ �      _newmode       __xi_a             �@ 8�         �@ Pw          �@ `�          A �          A 0^         A �K          HA p�      lA .debug_aranges .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges __mingw_invalidParameterHandler pre_c_init .rdata$.refptr.mingw_initltsdrot_force .rdata$.refptr.mingw_initltsdyn_force .rdata$.refptr.mingw_initltssuo_force .rdata$.refptr.mingw_initcharmax .rdata$.refptr.__image_base__ .rdata$.refptr.mingw_app_type managedapp .rdata$.refptr._fmode .rdata$.refptr._MINGW_INSTALL_DEBUG_MATHERR pre_cpp_init .rdata$.refptr._newmode startinfo .rdata$.refptr._dowildcard __tmainCRTStartu      p .rdata$.refptr.__native_startup_lock .rdata$.refptr.__native_startup_state has_cctor .rdata$.refptr.__dyn_tls_init_callback .rdata$.refptr.__mingw_oldexcpt_handler .rdata$.refptr.__imp___initenv .rdata$.refptr.__xc_z .rdata$.refptr.__xc_a .rdata$.refptr.__xi_z .rdata$.refptr.__xi_a WinMainCRTStartup .l_startw mainCRTStartup .rdata$.refptr._gnu_exception_handler .rdata$.refptr._matherr .CRT$XCAA .CRT$XIAA __gcc_register_frame __gcc_deregister_frame _ZStL19piecewise_construct _ZStL8__ioinit .rdata$.refptr._ZSt4cout .rdata$.refptr._ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_main .debug_info .debug_abbrev .debug_aranges .debug_line .debug_str .rdata$zzz .debug_frame _GLOBAL__sub_I_disk.cpp .data$_ZN14__gnu_internal9buf_wcerrE .data$_ZN14__gnu_internal8buf_wcinE .data$_ZN14__gnu_internal9buf_wcoutE .data$_ZN14__gnu_internal14buf_wcerr_syncE .data$_ZN14__gnu_internal13buf_wcin_syncE .data$_ZN14__gnu_internal14buf_wcout_syncE .da      ta$_ZN14__gnu_internal8buf_cerrE .data$_ZN14__gnu_internal7buf_cinE .data$_ZN14__gnu_internal8buf_coutE .data$_ZN14__gnu_internal13buf_cerr_syncE .data$_ZN14__gnu_internal12buf_cin_syncE .data$_ZN14__gnu_internal13buf_cout_syncE .data$_ZSt5wclog .data$_ZSt5wcerr .data$_ZSt5wcout .data$_ZSt4wcin .data$_ZSt4clog .data$_ZSt4cerr .data$_ZSt4cout .data$_ZSt3cin _ZNSt8ios_base4InitC2Ev .rdata$.refptr._ZNSt8ios_base4Init11_S_refcountE .rdata$.refptr._ZNSt8ios_base4Init20_S_synced_with_stdioE .rdata$.refptr._ZN14__gnu_internal13buf_cout_syncE .rdata$.refptr._ZTVSt15basic_streambufIcSt11char_traitsIcEE .rdata$.refptr._ZTVN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE .rdata$.refptr._ZN14__gnu_internal12buf_cin_syncE .rdata$.refptr._ZN14__gnu_internal13buf_cerr_syncE .rdata$.refptr._ZTVSo .rdata$.refptr._ZSt3cin .rdata$.refptr._ZTVSi .rdata$.refptr._ZSt4cerr .rdata$.refptr._ZSt4clog .rdata$.refptr._ZN14__gnu_internal14buf_wcout_syncE .rdata$.refptr._ZTVSt15basic_streambufIwSt11char_traitsIwEE .rdata$.ref      ptr._ZTVN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE .rdata$.refptr._ZN14__gnu_internal13buf_wcin_syncE .rdata$.refptr._ZN14__gnu_internal14buf_wcerr_syncE .rdata$.refptr._ZSt5wcout .rdata$.refptr._ZTVSt13basic_ostreamIwSt11char_traitsIwEE .rdata$.refptr._ZSt4wcin .rdata$.refptr._ZTVSt13basic_istreamIwSt11char_traitsIwEE .rdata$.refptr._ZSt5wcerr .rdata$.refptr._ZSt5wclog .rdata$.refptr._ZTVSt9basic_iosIcSt11char_traitsIcEE .rdata$.refptr._ZTVSt9basic_iosIwSt11char_traitsIwEE _ZNSt8ios_base4InitC1Ev _ZNSt8ios_base4InitD2Ev _ZNSt8ios_base4InitD1Ev _ZNSt8ios_base15sync_with_stdioEb .rdata$.refptr._ZN14__gnu_internal8buf_coutE .rdata$.refptr._ZN14__gnu_internal7buf_cinE .rdata$.refptr._ZN14__gnu_internal8buf_cerrE .rdata$.refptr._ZN14__gnu_internal9buf_wcoutE .rdata$.refptr._ZN14__gnu_internal8buf_wcinE .rdata$.refptr._ZN14__gnu_internal9buf_wcerrE .text$_ZNSt8ios_base4InitC2Ev .xdata$_ZNSt8ios_base4InitC2Ev .pdata$_ZNSt8ios_base4InitC2Ev .text$_ZNSt8ios_base4InitD2Ev .xdata$_ZNSt8ios_base4InitD      2Ev .pdata$_ZNSt8ios_base4InitD2Ev .text$_ZNSt8ios_base15sync_with_stdioEb .xdata$_ZNSt8ios_base15sync_with_stdioEb .pdata$_ZNSt8ios_base15sync_with_stdioEb .text$_ZNK9__gnu_cxx24__concurrence_lock_error4whatEv _ZNK9__gnu_cxx24__concurrence_lock_error4whatEv .text$_ZNK9__gnu_cxx26__concurrence_unlock_error4whatEv _ZNK9__gnu_cxx26__concurrence_unlock_error4whatEv _ZNSt6locale5facetD2Ev _ZNSt6locale5facetD1Ev _ZNSt6locale5facetD0Ev _ZNSt6locale5facet18_S_initialize_onceEv _ZZN12_GLOBAL__N_122get_locale_cache_mutexEvE18locale_cache_mutex .text$_ZN9__gnu_cxx24__concurrence_lock_errorD1Ev _ZN9__gnu_cxx24__concurrence_lock_errorD1Ev .rdata$_ZTVN9__gnu_cxx24__concurrence_lock_errorE .text$_ZN9__gnu_cxx24__concurrence_lock_errorD0Ev _ZN9__gnu_cxx24__concurrence_lock_errorD0Ev .text$_ZN9__gnu_cxx26__concurrence_unlock_errorD1Ev _ZN9__gnu_cxx26__concurrence_unlock_errorD1Ev .rdata$_ZTVN9__gnu_cxx26__concurrence_unlock_errorE .text$_ZN9__gnu_cxx26__concurrence_unlock_errorD0Ev _ZN9__gnu_cxx26__concurrence_unlock      _errorD0Ev .text$_ZN9__gnu_cxx13__scoped_lockD1Ev _ZN9__gnu_cxx13__scoped_lockD1Ev .rdata$_ZTIN9__gnu_cxx26__concurrence_unlock_errorE _ZNSt6localeC2ERKS_ _ZNSt6localeC1ERKS_ _ZNSt6localeC2EPNS_5_ImplE _ZNSt6localeC1EPNS_5_ImplE _ZNKSt6locale4nameB5cxx11Ev .rdata$.refptr._ZNSt6locale13_S_categoriesE _ZNKSt6localeeqERKS_ _ZNSt6locale21_S_normalize_categoryEi CSWTCH.42 _ZNSt6locale5facet15_S_get_c_localeEv _ZNSt6locale5facet13_S_get_c_nameEv _ZNSt6locale5_ImplD2Ev _ZNSt6locale5_ImplD1Ev _ZNSt6localeaSERKS_ _ZNSt6localeD2Ev _ZNSt6localeD1Ev _ZNSt6locale5_ImplC2ERKS0_y _ZNSt6locale5_ImplC1ERKS0_y _ZNKSt6locale2id5_M_idEv _ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE .rdata$.refptr._ZNSt6locale17_S_twinned_facetsE _ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE _ZNSt6locale5_Impl19_M_replace_categoryEPKS0_PKPKNS_2idE _ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEy _ZGVZN12_GLOBAL__N_122get_locale_cache_mutexEvE18locale_cache_mutex .rdata$_ZTIN9__gnu_cxx24__concurrence_lock_errorE .rdata      $_ZTSSt9exception .rdata$_ZTISt9exception .rdata$_ZTSNSt6locale5facetE .rdata$_ZTINSt6locale5facetE .rdata$_ZTSN9__gnu_cxx24__concurrence_lock_errorE .rdata$_ZTSN9__gnu_cxx26__concurrence_unlock_errorE .rdata$_ZTVNSt6locale5facetE .xdata$_ZNK9__gnu_cxx24__concurrence_lock_error4whatEv .pdata$_ZNK9__gnu_cxx24__concurrence_lock_error4whatEv .xdata$_ZNK9__gnu_cxx26__concurrence_unlock_error4whatEv .pdata$_ZNK9__gnu_cxx26__concurrence_unlock_error4whatEv .text$_ZNSt6locale5facetD2Ev .xdata$_ZNSt6locale5facetD2Ev .pdata$_ZNSt6locale5facetD2Ev .text$_ZNSt6locale5facetD0Ev .xdata$_ZNSt6locale5facetD0Ev .pdata$_ZNSt6locale5facetD0Ev .text$_ZNSt6locale5facet18_S_initialize_onceEv .xdata$_ZNSt6locale5facet18_S_initialize_onceEv .pdata$_ZNSt6locale5facet18_S_initialize_onceEv .text$__tcf_0 .xdata$__tcf_0 .pdata$__tcf_0 .xdata$_ZN9__gnu_cxx24__concurrence_lock_errorD1Ev .pdata$_ZN9__gnu_cxx24__concurrence_lock_errorD1Ev .xdata$_ZN9__gnu_cxx24__concurrence_lock_errorD0Ev .pdata$_ZN9__gnu_cxx24__concurrence_lock_er       rorD0Ev .xdata$_ZN9__gnu_cxx26__concurrence_unlock_errorD1Ev .pdata$_ZN9__gnu_cxx26__concurrence_unlock_errorD1Ev .xdata$_ZN9__gnu_cxx26__concurrence_unlock_errorD0Ev .pdata$_ZN9__gnu_cxx26__concurrence_unlock_errorD0Ev .xdata$_ZN9__gnu_cxx13__scoped_lockD1Ev .pdata$_ZN9__gnu_cxx13__scoped_lockD1Ev .text$_ZNSt6localeC2ERKS_ .xdata$_ZNSt6localeC2ERKS_ .pdata$_ZNSt6localeC2ERKS_ .text$_ZNSt6localeC2EPNS_5_ImplE .xdata$_ZNSt6localeC2EPNS_5_ImplE .pdata$_ZNSt6localeC2EPNS_5_ImplE .text$_ZNKSt6locale4nameB5cxx11Ev .xdata$_ZNKSt6locale4nameB5cxx11Ev .pdata$_ZNKSt6locale4nameB5cxx11Ev .text$_ZNKSt6localeeqERKS_ .xdata$_ZNKSt6localeeqERKS_ .pdata$_ZNKSt6localeeqERKS_ .text$_ZNSt6locale21_S_normalize_categoryEi .xdata$_ZNSt6locale21_S_normalize_categoryEi .pdata$_ZNSt6locale21_S_normalize_categoryEi .text$_ZNSt6locale5facet15_S_get_c_localeEv .xdata$_ZNSt6locale5facet15_S_get_c_localeEv .pdata$_ZNSt6locale5facet15_S_get_c_localeEv .text$_ZNSt6locale5facet13_S_get_c_nameEv .xdata$_ZNSt6locale5facet13_S_get_c_na!      meEv .pdata$_ZNSt6locale5facet13_S_get_c_nameEv .text$_ZNSt6locale5_ImplD2Ev .xdata$_ZNSt6locale5_ImplD2Ev .pdata$_ZNSt6locale5_ImplD2Ev .text$_ZNSt6localeaSERKS_ .xdata$_ZNSt6localeaSERKS_ .pdata$_ZNSt6localeaSERKS_ .text$_ZNSt6localeD2Ev .xdata$_ZNSt6localeD2Ev .pdata$_ZNSt6localeD2Ev .text$_ZNSt6locale5_ImplC2ERKS0_y .xdata$_ZNSt6locale5_ImplC2ERKS0_y .pdata$_ZNSt6locale5_ImplC2ERKS0_y .text$_ZNKSt6locale2id5_M_idEv .xdata$_ZNKSt6locale2id5_M_idEv .pdata$_ZNKSt6locale2id5_M_idEv .text$_ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE .xdata$_ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE .pdata$_ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE .text$_ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE .xdata$_ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE .pdata$_ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE .text$_ZNSt6locale5_Impl19_M_replace_categoryEPKS0_PKPKNS_2idE .xdata$_ZNSt6locale5_Impl19_M_replace_categoryEPKS0_PKPKNS_2idE .pdata$_ZNSt6locale5_Impl19_M"      _replace_categoryEPKS0_PKPKNS_2idE .text$_ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEy .xdata$_ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEy .pdata$_ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEy .rdata$CSWTCH.42 .data$_ZNSt6locale2id11_S_refcountE .data$_ZNSt6locale5facet7_S_onceE .rdata$_ZNSt6locale5facet9_S_c_nameE .data$_ZNSt6locale5facet11_S_c_localeE .data$_ZNSt6locale7_S_onceE .data$_ZNSt6locale9_S_globalE .data$_ZNSt6locale10_S_classicE .rdata$_ZNSt6locale3allE .rdata$_ZNSt6locale8messagesE .rdata$_ZNSt6locale8monetaryE .rdata$_ZNSt6locale4timeE .rdata$_ZNSt6locale7collateE .rdata$_ZNSt6locale7numericE .rdata$_ZNSt6locale5ctypeE .rdata$_ZNSt6locale4noneE .data$_ZGVZN12_GLOBAL__N_122get_locale_cache_mutexEvE18locale_cache_mutex .data$_ZZN12_GLOBAL__N_122get_locale_cache_mutexEvE18locale_cache_mutex _ZZN12_GLOBAL__N_116get_locale_mutexEvE12locale_mutex _ZN12_GLOBAL__N_116get_locale_mutexEv _ZGVZN12_GLOBAL__N_116get_locale_mutexEvE12locale_mutex .text$_ZN9__gnu_cxx30__throw_concurrenc#      e_lock_errorEv _ZN9__gnu_cxx30__throw_concurrence_lock_errorEv _ZNSt6locale5_ImplC2Ey _ZN12_GLOBAL__N_19facet_vecE _ZN12_GLOBAL__N_19cache_vecE _ZN12_GLOBAL__N_18name_vecE _ZN12_GLOBAL__N_16name_cE _ZN12_GLOBAL__N_17ctype_cE .rdata$.refptr._ZNSt5ctypeIcE2idE _ZN12_GLOBAL__N_19codecvt_cE .rdata$.refptr._ZNSt7codecvtIcciE2idE .rdata$.refptr._ZTVSt16__numpunct_cacheIcE _ZN12_GLOBAL__N_116numpunct_cache_cE _ZN12_GLOBAL__N_110numpunct_cE .rdata$.refptr._ZTVNSt7__cxx118numpunctIcEE .rdata$.refptr._ZNSt7__cxx118numpunctIcE2idE .rdata$.refptr._ZTVSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZN12_GLOBAL__N_19num_get_cE .rdata$.refptr._ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZN12_GLOBAL__N_19num_put_cE .rdata$.refptr._ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVNSt7__cxx117collateIcEE _ZN12_GLOBAL__N_19collate_cE .rdata$.refptr._ZNSt7__cxx117collateIcE2idE .r$      data$.refptr._ZTVSt18__moneypunct_cacheIcLb0EE _ZN12_GLOBAL__N_119moneypunct_cache_cfE _ZN12_GLOBAL__N_113moneypunct_cfE .rdata$.refptr._ZTVNSt7__cxx1110moneypunctIcLb0EEE .rdata$.refptr._ZNSt7__cxx1110moneypunctIcLb0EE2idE .rdata$.refptr._ZTVSt18__moneypunct_cacheIcLb1EE _ZN12_GLOBAL__N_119moneypunct_cache_ctE _ZN12_GLOBAL__N_113moneypunct_ctE .rdata$.refptr._ZTVNSt7__cxx1110moneypunctIcLb1EEE .rdata$.refptr._ZNSt7__cxx1110moneypunctIcLb1EE2idE .rdata$.refptr._ZTVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZN12_GLOBAL__N_111money_get_cE .rdata$.refptr._ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE _ZN12_GLOBAL__N_111money_put_cE .rdata$.refptr._ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVSt17__timepunct_cacheIcE _ZN12_GLOBAL__N_117timepunct_cache_cE _ZN12_GLOBAL__N_111timepunct_cE .rdata$.refptr._ZNSt11__timepu%      nctIcE2idE .rdata$.refptr._ZTVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZN12_GLOBAL__N_110time_get_cE .rdata$.refptr._ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZN12_GLOBAL__N_110time_put_cE .rdata$.refptr._ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZN12_GLOBAL__N_110messages_cE .rdata$.refptr._ZNSt7__cxx118messagesIcE2idE _ZN12_GLOBAL__N_17ctype_wE .rdata$.refptr._ZNSt5ctypeIwE2idE _ZN12_GLOBAL__N_19codecvt_wE .rdata$.refptr._ZNSt7codecvtIwciE2idE .rdata$.refptr._ZTVSt16__numpunct_cacheIwE _ZN12_GLOBAL__N_116numpunct_cache_wE _ZN12_GLOBAL__N_110numpunct_wE .rdata$.refptr._ZTVNSt7__cxx118numpunctIwEE .rdata$.refptr._ZNSt7__cxx118numpunctIwE2idE .rdata$.refptr._ZTVSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZN12_GLOBAL__N_19num_get_wE .rdata$.refptr._ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._Z&      TVSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZN12_GLOBAL__N_19num_put_wE .rdata$.refptr._ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._ZTVNSt7__cxx117collateIwEE _ZN12_GLOBAL__N_19collate_wE .rdata$.refptr._ZNSt7__cxx117collateIwE2idE .rdata$.refptr._ZTVSt18__moneypunct_cacheIwLb0EE _ZN12_GLOBAL__N_119moneypunct_cache_wfE _ZN12_GLOBAL__N_113moneypunct_wfE .rdata$.refptr._ZTVNSt7__cxx1110moneypunctIwLb0EEE .rdata$.refptr._ZNSt7__cxx1110moneypunctIwLb0EE2idE .rdata$.refptr._ZTVSt18__moneypunct_cacheIwLb1EE _ZN12_GLOBAL__N_119moneypunct_cache_wtE _ZN12_GLOBAL__N_113moneypunct_wtE .rdata$.refptr._ZTVNSt7__cxx1110moneypunctIwLb1EEE .rdata$.refptr._ZNSt7__cxx1110moneypunctIwLb1EE2idE .rdata$.refptr._ZTVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZN12_GLOBAL__N_111money_get_wE .rdata$.refptr._ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._ZTVNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwS'      t11char_traitsIwEEEE _ZN12_GLOBAL__N_111money_put_wE .rdata$.refptr._ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._ZTVSt17__timepunct_cacheIwE _ZN12_GLOBAL__N_117timepunct_cache_wE _ZN12_GLOBAL__N_111timepunct_wE .rdata$.refptr._ZNSt11__timepunctIwE2idE .rdata$.refptr._ZTVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZN12_GLOBAL__N_110time_get_wE .rdata$.refptr._ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._ZTVSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZN12_GLOBAL__N_110time_put_wE .rdata$.refptr._ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZN12_GLOBAL__N_110messages_wE .rdata$.refptr._ZNSt7__cxx118messagesIwE2idE .rdata$.refptr._ZTVSt7codecvtIDsciE _ZN12_GLOBAL__N_111codecvt_c16E .rdata$.refptr._ZNSt7codecvtIDsciE2idE .rdata$.refptr._ZTVSt7codecvtIDiciE _ZN12_GLOBAL__N_111codecvt_c32E .rdata$.refptr._ZNSt7codecvtIDiciE2idE _ZNSt6locale5_ImplC1Ey _ZNSt6l(      ocale18_S_initialize_onceEv _ZN12_GLOBAL__N_113c_locale_implE .rdata$.refptr._ZNSt6locale10_S_classicE .rdata$.refptr._ZNSt6locale9_S_globalE _ZNSt6locale13_S_initializeEv .rdata$.refptr._ZNSt6locale7_S_onceE _ZNSt6localeC2Ev _ZNSt6localeC1Ev _ZNSt6locale7classicEv _ZN12_GLOBAL__N_18c_localeE _ZNSt6locale6globalERKS_ .text$_ZN12_GLOBAL__N_116get_locale_mutexEv .xdata$_ZN12_GLOBAL__N_116get_locale_mutexEv .pdata$_ZN12_GLOBAL__N_116get_locale_mutexEv .xdata$_ZN9__gnu_cxx30__throw_concurrence_lock_errorEv .pdata$_ZN9__gnu_cxx30__throw_concurrence_lock_errorEv .text$_ZNSt6locale5_ImplC2Ey .xdata$_ZNSt6locale5_ImplC2Ey .pdata$_ZNSt6locale5_ImplC2Ey .text$_ZNSt6locale18_S_initialize_onceEv .xdata$_ZNSt6locale18_S_initialize_onceEv .pdata$_ZNSt6locale18_S_initialize_onceEv .text$_ZNSt6locale13_S_initializeEv .xdata$_ZNSt6locale13_S_initializeEv .pdata$_ZNSt6locale13_S_initializeEv .text$_ZNSt6localeC2Ev .xdata$_ZNSt6localeC2Ev .pdata$_ZNSt6localeC2Ev .text$_ZNSt6locale7classicEv .xdata$_ZNSt6locale7classicEv)       .pdata$_ZNSt6locale7classicEv .text$_ZNSt6locale6globalERKS_ .xdata$_ZNSt6locale6globalERKS_ .pdata$_ZNSt6locale6globalERKS_ .rdata$_ZNSt6locale17_S_twinned_facetsE .rdata$_ZNSt6locale5_Impl19_S_facet_categoriesE .rdata$_ZNSt6locale5_Impl14_S_id_messagesE .rdata$_ZNSt6locale5_Impl14_S_id_monetaryE .rdata$_ZNSt6locale5_Impl10_S_id_timeE .rdata$_ZNSt6locale5_Impl13_S_id_collateE .rdata$_ZNSt6locale5_Impl13_S_id_numericE .rdata$_ZNSt6locale5_Impl11_S_id_ctypeE .data$_ZN12_GLOBAL__N_117timepunct_cache_wE .data$_ZN12_GLOBAL__N_119moneypunct_cache_wfE .data$_ZN12_GLOBAL__N_119moneypunct_cache_wtE .data$_ZN12_GLOBAL__N_116numpunct_cache_wE .data$_ZN12_GLOBAL__N_117timepunct_cache_cE .data$_ZN12_GLOBAL__N_119moneypunct_cache_cfE .data$_ZN12_GLOBAL__N_119moneypunct_cache_ctE .data$_ZN12_GLOBAL__N_116numpunct_cache_cE .data$_ZN12_GLOBAL__N_111codecvt_c32E .data$_ZN12_GLOBAL__N_111codecvt_c16E .data$_ZN12_GLOBAL__N_110messages_wE .data$_ZN12_GLOBAL__N_110time_put_wE .data$_ZN12_GLOBAL__N_110time_get_wE .data$_Z*      N12_GLOBAL__N_111timepunct_wE .data$_ZN12_GLOBAL__N_111money_put_wE .data$_ZN12_GLOBAL__N_111money_get_wE .data$_ZN12_GLOBAL__N_113moneypunct_wfE .data$_ZN12_GLOBAL__N_113moneypunct_wtE .data$_ZN12_GLOBAL__N_19codecvt_wE .data$_ZN12_GLOBAL__N_19num_put_wE .data$_ZN12_GLOBAL__N_19num_get_wE .data$_ZN12_GLOBAL__N_110numpunct_wE .data$_ZN12_GLOBAL__N_19collate_wE .data$_ZN12_GLOBAL__N_17ctype_wE .data$_ZN12_GLOBAL__N_110messages_cE .data$_ZN12_GLOBAL__N_110time_put_cE .data$_ZN12_GLOBAL__N_110time_get_cE .data$_ZN12_GLOBAL__N_111timepunct_cE .data$_ZN12_GLOBAL__N_111money_put_cE .data$_ZN12_GLOBAL__N_111money_get_cE .data$_ZN12_GLOBAL__N_113moneypunct_cfE .data$_ZN12_GLOBAL__N_113moneypunct_ctE .data$_ZN12_GLOBAL__N_19codecvt_cE .data$_ZN12_GLOBAL__N_19num_put_cE .data$_ZN12_GLOBAL__N_19num_get_cE .data$_ZN12_GLOBAL__N_110numpunct_cE .data$_ZN12_GLOBAL__N_19collate_cE .data$_ZN12_GLOBAL__N_17ctype_cE .data$_ZN12_GLOBAL__N_19cache_vecE .data$_ZN12_GLOBAL__N_19facet_vecE .data$_ZN12_GLOBAL__N_16name_cE .da+      ta$_ZN12_GLOBAL__N_18name_vecE .data$_ZN12_GLOBAL__N_18c_localeE .data$_ZN12_GLOBAL__N_113c_locale_implE .data$_ZGVZN12_GLOBAL__N_116get_locale_mutexEvE12locale_mutex .data$_ZZN12_GLOBAL__N_116get_locale_mutexEvE12locale_mutex _ZNSt7__cxx1110moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .rdata$.refptr._ZNSt10money_base18_S_default_patternE .rdata$.refptr._ZNSt10money_base8_S_atomsE _ZNSt7__cxx1110moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc _ZNSt7__cxx1110moneypunctIcLb1EED2Ev _ZNSt7__cxx1110moneypunctIcLb1EED1Ev _ZNSt7__cxx1110moneypunctIcLb1EED0Ev _ZNSt7__cxx1110moneypunctIcLb0EED2Ev _ZNSt7__cxx1110moneypunctIcLb0EED1Ev _ZNSt7__cxx1110moneypunctIcLb0EED0Ev _ZNSt7__cxx1110moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc _ZNSt7__cxx1110moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc _ZNSt7__cxx1110moneypunctIwLb1EED2Ev _ZNSt7__cxx1110moneypunctIwLb1EED1Ev _ZNSt7__cxx1110moneypunctIwLb1EED0Ev _ZNSt7__cxx1110moneypunctIwLb0EED2Ev _ZNSt7__cxx1110moneypunctIwLb0EED1Ev _ZNSt7__cxx1110moneypunct,      IwLb0EED0Ev .text$_ZNSt7__cxx1110moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt7__cxx1110moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt7__cxx1110moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt7__cxx1110moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt7__cxx1110moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt7__cxx1110moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt7__cxx1110moneypunctIcLb1EED2Ev .xdata$_ZNSt7__cxx1110moneypunctIcLb1EED2Ev .pdata$_ZNSt7__cxx1110moneypunctIcLb1EED2Ev .text$_ZNSt7__cxx1110moneypunctIcLb1EED0Ev .xdata$_ZNSt7__cxx1110moneypunctIcLb1EED0Ev .pdata$_ZNSt7__cxx1110moneypunctIcLb1EED0Ev .text$_ZNSt7__cxx1110moneypunctIcLb0EED2Ev .xdata$_ZNSt7__cxx1110moneypunctIcLb0EED2Ev .pdata$_ZNSt7__cxx1110moneypunctIcLb0EED2Ev .text$_ZNSt7__cxx1110moneypunctIcLb0EED0Ev .xdata$_ZNSt7__cxx1110moneypunctIcLb0EED0Ev .pdata$_ZNSt7__cxx1110moneypunctIcLb0EED0Ev .text$_ZNSt7__cxx1110moneypunctIwLb1EE24_M_initial-      ize_moneypunctEPiPKc .xdata$_ZNSt7__cxx1110moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt7__cxx1110moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt7__cxx1110moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt7__cxx1110moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt7__cxx1110moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt7__cxx1110moneypunctIwLb1EED2Ev .xdata$_ZNSt7__cxx1110moneypunctIwLb1EED2Ev .pdata$_ZNSt7__cxx1110moneypunctIwLb1EED2Ev .text$_ZNSt7__cxx1110moneypunctIwLb1EED0Ev .xdata$_ZNSt7__cxx1110moneypunctIwLb1EED0Ev .pdata$_ZNSt7__cxx1110moneypunctIwLb1EED0Ev .text$_ZNSt7__cxx1110moneypunctIwLb0EED2Ev .xdata$_ZNSt7__cxx1110moneypunctIwLb0EED2Ev .pdata$_ZNSt7__cxx1110moneypunctIwLb0EED2Ev .text$_ZNSt7__cxx1110moneypunctIwLb0EED0Ev .xdata$_ZNSt7__cxx1110moneypunctIwLb0EED0Ev .pdata$_ZNSt7__cxx1110moneypunctIwLb0EED0Ev .text$_ZNSt18__moneypunct_cacheIcLb1EED1Ev _ZNSt18__moneypunct_cacheIcLb1EED1Ev .rdata$_ZTVSt18__moneypunct_cach.      eIcLb1EE .text$_ZNSt18__moneypunct_cacheIcLb1EED0Ev _ZNSt18__moneypunct_cacheIcLb1EED0Ev .text$_ZNSt18__moneypunct_cacheIcLb0EED1Ev _ZNSt18__moneypunct_cacheIcLb0EED1Ev .rdata$_ZTVSt18__moneypunct_cacheIcLb0EE .text$_ZNSt18__moneypunct_cacheIcLb0EED0Ev _ZNSt18__moneypunct_cacheIcLb0EED0Ev .text$_ZNSt18__moneypunct_cacheIwLb1EED1Ev _ZNSt18__moneypunct_cacheIwLb1EED1Ev .rdata$_ZTVSt18__moneypunct_cacheIwLb1EE .text$_ZNSt18__moneypunct_cacheIwLb1EED0Ev _ZNSt18__moneypunct_cacheIwLb1EED0Ev .text$_ZNSt18__moneypunct_cacheIwLb0EED1Ev _ZNSt18__moneypunct_cacheIwLb0EED1Ev .rdata$_ZTVSt18__moneypunct_cacheIwLb0EE .text$_ZNSt18__moneypunct_cacheIwLb0EED0Ev _ZNSt18__moneypunct_cacheIwLb0EED0Ev _ZNSt10money_base20_S_construct_patternEccc _ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc _ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc _ZNSt10moneypunctIcLb1EED2Ev .rdata$.refptr._ZTVSt10moneypunctIcLb1EE _ZNSt10moneypunctIcLb1EED1Ev _ZNSt10moneypunctIcLb1EED0Ev _ZNSt10moneypunctIcLb0EED2Ev .rdata$.r/      efptr._ZTVSt10moneypunctIcLb0EE _ZNSt10moneypunctIcLb0EED1Ev _ZNSt10moneypunctIcLb0EED0Ev _ZNSt10moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc _ZNSt10moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc _ZNSt10moneypunctIwLb1EED2Ev .rdata$.refptr._ZTVSt10moneypunctIwLb1EE _ZNSt10moneypunctIwLb1EED1Ev _ZNSt10moneypunctIwLb1EED0Ev _ZNSt10moneypunctIwLb0EED2Ev .rdata$.refptr._ZTVSt10moneypunctIwLb0EE _ZNSt10moneypunctIwLb0EED1Ev _ZNSt10moneypunctIwLb0EED0Ev .rdata$_ZTSSt18__moneypunct_cacheIcLb1EE .rdata$_ZTISt18__moneypunct_cacheIcLb1EE .rdata$_ZTSSt18__moneypunct_cacheIcLb0EE .rdata$_ZTISt18__moneypunct_cacheIcLb0EE .rdata$_ZTSSt18__moneypunct_cacheIwLb1EE .rdata$_ZTISt18__moneypunct_cacheIwLb1EE .rdata$_ZTSSt18__moneypunct_cacheIwLb0EE .rdata$_ZTISt18__moneypunct_cacheIwLb0EE .xdata$_ZNSt18__moneypunct_cacheIcLb1EED1Ev .pdata$_ZNSt18__moneypunct_cacheIcLb1EED1Ev .xdata$_ZNSt18__moneypunct_cacheIcLb1EED0Ev .pdata$_ZNSt18__moneypunct_cacheIcLb1EED0Ev .xdata$_ZNSt18__moneypunct_cacheIcLb0EED1Ev .pdata$_0      ZNSt18__moneypunct_cacheIcLb0EED1Ev .xdata$_ZNSt18__moneypunct_cacheIcLb0EED0Ev .pdata$_ZNSt18__moneypunct_cacheIcLb0EED0Ev .xdata$_ZNSt18__moneypunct_cacheIwLb1EED1Ev .pdata$_ZNSt18__moneypunct_cacheIwLb1EED1Ev .xdata$_ZNSt18__moneypunct_cacheIwLb1EED0Ev .pdata$_ZNSt18__moneypunct_cacheIwLb1EED0Ev .xdata$_ZNSt18__moneypunct_cacheIwLb0EED1Ev .pdata$_ZNSt18__moneypunct_cacheIwLb0EED1Ev .xdata$_ZNSt18__moneypunct_cacheIwLb0EED0Ev .pdata$_ZNSt18__moneypunct_cacheIwLb0EED0Ev .text$_ZNSt10money_base20_S_construct_patternEccc .xdata$_ZNSt10money_base20_S_construct_patternEccc .pdata$_ZNSt10money_base20_S_construct_patternEccc .text$_ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc .text$1      _ZNSt10moneypunctIcLb1EED2Ev .xdata$_ZNSt10moneypunctIcLb1EED2Ev .pdata$_ZNSt10moneypunctIcLb1EED2Ev .text$_ZNSt10moneypunctIcLb1EED0Ev .xdata$_ZNSt10moneypunctIcLb1EED0Ev .pdata$_ZNSt10moneypunctIcLb1EED0Ev .text$_ZNSt10moneypunctIcLb0EED2Ev .xdata$_ZNSt10moneypunctIcLb0EED2Ev .pdata$_ZNSt10moneypunctIcLb0EED2Ev .text$_ZNSt10moneypunctIcLb0EED0Ev .xdata$_ZNSt10moneypunctIcLb0EED0Ev .pdata$_ZNSt10moneypunctIcLb0EED0Ev .text$_ZNSt10moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt10moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt10moneypunctIwLb1EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt10moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .xdata$_ZNSt10moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .pdata$_ZNSt10moneypunctIwLb0EE24_M_initialize_moneypunctEPiPKc .text$_ZNSt10moneypunctIwLb1EED2Ev .xdata$_ZNSt10moneypunctIwLb1EED2Ev .pdata$_ZNSt10moneypunctIwLb1EED2Ev .text$_ZNSt10moneypunctIwLb1EED0Ev .xdata$_ZNSt10moneypunctIwLb1EED0Ev .pdata$_ZNSt10moneypunctIwLb1EED0E2      v .text$_ZNSt10moneypunctIwLb0EED2Ev .xdata$_ZNSt10moneypunctIwLb0EED2Ev .pdata$_ZNSt10moneypunctIwLb0EED2Ev .text$_ZNSt10moneypunctIwLb0EED0Ev .xdata$_ZNSt10moneypunctIwLb0EED0Ev .pdata$_ZNSt10moneypunctIwLb0EED0Ev _ZNSt7__cxx118numpunctIcE22_M_initialize_numpunctEPi .rdata$.refptr._ZNSt10__num_base12_S_atoms_outE .rdata$.refptr._ZNSt10__num_base11_S_atoms_inE _ZNSt7__cxx118numpunctIcED2Ev _ZNSt7__cxx118numpunctIcED1Ev _ZNSt7__cxx118numpunctIcED0Ev _ZNSt7__cxx118numpunctIwE22_M_initialize_numpunctEPi _ZNSt7__cxx118numpunctIwED2Ev _ZNSt7__cxx118numpunctIwED1Ev _ZNSt7__cxx118numpunctIwED0Ev .text$_ZNSt7__cxx118numpunctIcE22_M_initialize_numpunctEPi .xdata$_ZNSt7__cxx118numpunctIcE22_M_initialize_numpunctEPi .pdata$_ZNSt7__cxx118numpunctIcE22_M_initialize_numpunctEPi .text$_ZNSt7__cxx118numpunctIcED2Ev .xdata$_ZNSt7__cxx118numpunctIcED2Ev .pdata$_ZNSt7__cxx118numpunctIcED2Ev .text$_ZNSt7__cxx118numpunctIcED0Ev .xdata$_ZNSt7__cxx118numpunctIcED0Ev .pdata$_ZNSt7__cxx118numpunctIcED0Ev .text$_ZNSt7__cxx1183      numpunctIwE22_M_initialize_numpunctEPi .xdata$_ZNSt7__cxx118numpunctIwE22_M_initialize_numpunctEPi .pdata$_ZNSt7__cxx118numpunctIwE22_M_initialize_numpunctEPi .text$_ZNSt7__cxx118numpunctIwED2Ev .xdata$_ZNSt7__cxx118numpunctIwED2Ev .pdata$_ZNSt7__cxx118numpunctIwED2Ev .text$_ZNSt7__cxx118numpunctIwED0Ev .xdata$_ZNSt7__cxx118numpunctIwED0Ev .pdata$_ZNSt7__cxx118numpunctIwED0Ev .text$_ZNSt16__numpunct_cacheIcED1Ev _ZNSt16__numpunct_cacheIcED1Ev .rdata$_ZTVSt16__numpunct_cacheIcE .text$_ZNSt16__numpunct_cacheIcED0Ev _ZNSt16__numpunct_cacheIcED0Ev .text$_ZNSt16__numpunct_cacheIwED1Ev _ZNSt16__numpunct_cacheIwED1Ev .rdata$_ZTVSt16__numpunct_cacheIwE .text$_ZNSt16__numpunct_cacheIwED0Ev _ZNSt16__numpunct_cacheIwED0Ev _ZNSt8numpunctIcE22_M_initialize_numpunctEPi _ZNSt8numpunctIcED2Ev .rdata$.refptr._ZTVSt8numpunctIcE _ZNSt8numpunctIcED1Ev _ZNSt8numpunctIcED0Ev _ZNSt8numpunctIwE22_M_initialize_numpunctEPi _ZNSt8numpunctIwED2Ev .rdata$.refptr._ZTVSt8numpunctIwE _ZNSt8numpunctIwED1Ev _ZNSt8numpunctIwED0Ev .rdat4      a$_ZTSSt16__numpunct_cacheIcE .rdata$_ZTISt16__numpunct_cacheIcE .rdata$_ZTSSt16__numpunct_cacheIwE .rdata$_ZTISt16__numpunct_cacheIwE .xdata$_ZNSt16__numpunct_cacheIcED1Ev .pdata$_ZNSt16__numpunct_cacheIcED1Ev .xdata$_ZNSt16__numpunct_cacheIcED0Ev .pdata$_ZNSt16__numpunct_cacheIcED0Ev .xdata$_ZNSt16__numpunct_cacheIwED1Ev .pdata$_ZNSt16__numpunct_cacheIwED1Ev .xdata$_ZNSt16__numpunct_cacheIwED0Ev .pdata$_ZNSt16__numpunct_cacheIwED0Ev .text$_ZNSt8numpunctIcE22_M_initialize_numpunctEPi .xdata$_ZNSt8numpunctIcE22_M_initialize_numpunctEPi .pdata$_ZNSt8numpunctIcE22_M_initialize_numpunctEPi .text$_ZNSt8numpunctIcED2Ev .xdata$_ZNSt8numpunctIcED2Ev .pdata$_ZNSt8numpunctIcED2Ev .text$_ZNSt8numpunctIcED0Ev .xdata$_ZNSt8numpunctIcED0Ev .pdata$_ZNSt8numpunctIcED0Ev .text$_ZNSt8numpunctIwE22_M_initialize_numpunctEPi .xdata$_ZNSt8numpunctIwE22_M_initialize_numpunctEPi .pdata$_ZNSt8numpunctIwE22_M_initialize_numpunctEPi .text$_ZNSt8numpunctIwED2Ev .xdata$_ZNSt8numpunctIwED2Ev .pdata$_ZNSt8numpunctIwED2Ev .text$_ZN5      St8numpunctIwED0Ev .xdata$_ZNSt8numpunctIwED0Ev .pdata$_ZNSt8numpunctIwED0Ev _ZNSt12_GLOBAL__N_120read_utf8_code_pointERNS_5rangeIKcLb1EEEm _ZNKSt7codecvtIDsciE10do_unshiftERiPcS2_RS2_ _ZNKSt25__codecvt_utf8_utf16_baseIwE10do_unshiftERiPcS2_RS2_ _ZNKSt20__codecvt_utf16_baseIwE10do_unshiftERiPcS2_RS2_ _ZNKSt19__codecvt_utf8_baseIwE10do_unshiftERiPcS2_RS2_ _ZNKSt25__codecvt_utf8_utf16_baseIDiE10do_unshiftERiPcS2_RS2_ _ZNKSt20__codecvt_utf16_baseIDiE10do_unshiftERiPcS2_RS2_ _ZNKSt19__codecvt_utf8_baseIDiE10do_unshiftERiPcS2_RS2_ _ZNKSt25__codecvt_utf8_utf16_baseIDsE10do_unshiftERiPcS2_RS2_ _ZNKSt20__codecvt_utf16_baseIDsE10do_unshiftERiPcS2_RS2_ _ZNKSt19__codecvt_utf8_baseIDsE10do_unshiftERiPcS2_RS2_ _ZNKSt7codecvtIDiciE10do_unshiftERiPcS2_RS2_ _ZNKSt7codecvtIDsciE11do_encodingEv _ZNKSt25__codecvt_utf8_utf16_baseIwE11do_encodingEv _ZNKSt20__codecvt_utf16_baseIwE11do_encodingEv _ZNKSt19__codecvt_utf8_baseIwE11do_encodingEv _ZNKSt25__codecvt_utf8_utf16_baseIDiE11do_encodingEv _ZNKSt20__codecvt_utf16_baseID6      iE11do_encodingEv _ZNKSt19__codecvt_utf8_baseIDiE11do_encodingEv _ZNKSt25__codecvt_utf8_utf16_baseIDsE11do_encodingEv _ZNKSt20__codecvt_utf16_baseIDsE11do_encodingEv _ZNKSt19__codecvt_utf8_baseIDsE11do_encodingEv _ZNKSt7codecvtIDiciE11do_encodingEv _ZNKSt7codecvtIDsciE16do_always_noconvEv _ZNKSt25__codecvt_utf8_utf16_baseIwE16do_always_noconvEv _ZNKSt20__codecvt_utf16_baseIwE16do_always_noconvEv _ZNKSt19__codecvt_utf8_baseIwE16do_always_noconvEv _ZNKSt25__codecvt_utf8_utf16_baseIDiE16do_always_noconvEv _ZNKSt20__codecvt_utf16_baseIDiE16do_always_noconvEv _ZNKSt19__codecvt_utf8_baseIDiE16do_always_noconvEv _ZNKSt25__codecvt_utf8_utf16_baseIDsE16do_always_noconvEv _ZNKSt20__codecvt_utf16_baseIDsE16do_always_noconvEv _ZNKSt19__codecvt_utf8_baseIDsE16do_always_noconvEv _ZNKSt7codecvtIDiciE16do_always_noconvEv _ZNKSt7codecvtIDsciE13do_max_lengthEv _ZNKSt7codecvtIDiciE13do_max_lengthEv _ZNKSt19__codecvt_utf8_baseIDsE13do_max_lengthEv _ZNKSt19__codecvt_utf8_baseIDiE13do_max_lengthEv _ZNKSt19__codecvt_utf8_ba7      seIwE13do_max_lengthEv _ZNKSt20__codecvt_utf16_baseIDsE13do_max_lengthEv _ZNKSt20__codecvt_utf16_baseIDiE13do_max_lengthEv _ZNKSt20__codecvt_utf16_baseIwE13do_max_lengthEv _ZNKSt25__codecvt_utf8_utf16_baseIDsE13do_max_lengthEv _ZNKSt25__codecvt_utf8_utf16_baseIDiE13do_max_lengthEv _ZNKSt25__codecvt_utf8_utf16_baseIwE13do_max_lengthEv _ZNSt7codecvtIDsciED2Ev .rdata$_ZTVSt23__codecvt_abstract_baseIDsciE _ZNSt7codecvtIDsciED1Ev _ZNSt19__codecvt_utf8_baseIDsED2Ev _ZNSt19__codecvt_utf8_baseIDsED1Ev _ZNSt20__codecvt_utf16_baseIDsED2Ev _ZNSt20__codecvt_utf16_baseIDsED1Ev _ZNSt25__codecvt_utf8_utf16_baseIDsED2Ev _ZNSt25__codecvt_utf8_utf16_baseIDsED1Ev _ZNSt7codecvtIDiciED2Ev .rdata$_ZTVSt23__codecvt_abstract_baseIDiciE _ZNSt7codecvtIDiciED1Ev _ZNSt19__codecvt_utf8_baseIDiED2Ev _ZNSt19__codecvt_utf8_baseIDiED1Ev _ZNSt20__codecvt_utf16_baseIDiED2Ev _ZNSt20__codecvt_utf16_baseIDiED1Ev _ZNSt25__codecvt_utf8_utf16_baseIDiED2Ev _ZNSt25__codecvt_utf8_utf16_baseIDiED1Ev _ZNSt7codecvtIDsciED0Ev _ZNSt19__codecvt_utf8_8      baseIDsED0Ev _ZNSt20__codecvt_utf16_baseIDsED0Ev _ZNSt25__codecvt_utf8_utf16_baseIDsED0Ev _ZNSt7codecvtIDiciED0Ev _ZNSt19__codecvt_utf8_baseIDiED0Ev _ZNSt20__codecvt_utf16_baseIDiED0Ev _ZNSt25__codecvt_utf8_utf16_baseIDiED0Ev _ZNSt12_GLOBAL__N_18read_bomIKDsLb0ELy2EEEbRNS_5rangeIT_XT0_EEERAT1__Kh _ZNSt12_GLOBAL__N_121read_utf16_code_pointILb0EEEDiRNS_5rangeIKDsXT_EEEmSt12codecvt_mode _ZNSt19__codecvt_utf8_baseIwED2Ev .rdata$_ZTVSt19__codecvt_utf8_baseIwE _ZNSt19__codecvt_utf8_baseIwED1Ev _ZNSt19__codecvt_utf8_baseIwED0Ev _ZNSt20__codecvt_utf16_baseIwED2Ev .rdata$_ZTVSt20__codecvt_utf16_baseIwE _ZNSt20__codecvt_utf16_baseIwED1Ev _ZNSt20__codecvt_utf16_baseIwED0Ev _ZNSt25__codecvt_utf8_utf16_baseIwED2Ev .rdata$_ZTVSt25__codecvt_utf8_utf16_baseIwE _ZNSt25__codecvt_utf8_utf16_baseIwED1Ev _ZNSt25__codecvt_utf8_utf16_baseIwED0Ev _ZNSt12_GLOBAL__N_121write_utf8_code_pointERNS_5rangeIcLb1EEEDi _ZNSt12_GLOBAL__N_115write_utf16_bomILb0EEEbRNS_5rangeIDsXT_EEESt12codecvt_mode _ZNSt12_GLOBAL__N_1L11utf16le_bomE _Z9      NSt12_GLOBAL__N_1L9utf16_bomE _ZNKSt20__codecvt_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ _ZNSt12_GLOBAL__N_114write_utf8_bomERNS_5rangeIcLb1EEESt12codecvt_mode.part.19 _ZNSt12_GLOBAL__N_1L8utf8_bomE _ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE.part.20 _ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE _ZNKSt25__codecvt_utf8_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ _ZNKSt19__codecvt_utf8_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ _ZNKSt19__codecvt_utf8_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ _ZNKSt7codecvtIDsciE6do_outERiPKDsS3_RS3_PcS5_RS5_ _ZNKSt19__codecvt_utf8_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ _ZNSt12_GLOBAL__N_114read_utf16_bomILb0EEEvRNS_5rangeIKDsXT_EEERSt12codecvt_mode _ZNKSt20__codecvt_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ _ZNKSt20__codecvt_utf16_baseIDiE9do_lengthERiPKcS3_y _ZNSt12_GLOBAL__N_17ucs2_inERNS_5rangeIKDsLb0EEERNS0_I:      DsLb1EEEDiSt12codecvt_mode _ZNKSt20__codecvt_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ _ZNKSt20__codecvt_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ _ZNSt12_GLOBAL__N_19ucs2_spanERNS_5rangeIKDsLb0EEEyDiSt12codecvt_mode _ZNKSt20__codecvt_utf16_baseIDsE9do_lengthERiPKcS3_y _ZNKSt20__codecvt_utf16_baseIwE9do_lengthERiPKcS3_y _ZNSt12_GLOBAL__N_18ucs2_outERNS_5rangeIKDsLb1EEERNS0_IDsLb0EEEDiSt12codecvt_mode.part.23 _ZNKSt20__codecvt_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ _ZNKSt25__codecvt_utf8_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ _ZNKSt25__codecvt_utf8_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ _ZNSt12_GLOBAL__N_18read_bomIKcLb1ELy3EEEbRNS_5rangeIT_XT0_EEERAT1__Kh.constprop.29 _ZNKSt25__codecvt_utf8_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ _ZNKSt25__codecvt_utf8_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ _ZNSt12_GLOBAL__N_19ucs2_spanEPKcS1_yDiSt12codecvt_mode _ZNKSt19__codecvt_utf8_baseIDsE9do_lengthERiPKcS3_y _ZNKSt19__codecvt_utf8_baseIwE9do_lengthERiPKcS3_y _ZNSt12_GLOBAL__N_110utf16_spa;      nEPKcS1_yDiSt12codecvt_mode _ZNKSt7codecvtIDsciE9do_lengthERiPKcS3_y _ZNKSt25__codecvt_utf8_utf16_baseIDsE9do_lengthERiPKcS3_y _ZNKSt25__codecvt_utf8_utf16_baseIDiE9do_lengthERiPKcS3_y _ZNKSt25__codecvt_utf8_utf16_baseIwE9do_lengthERiPKcS3_y _ZNSt12_GLOBAL__N_18utf16_inIDsEENSt12codecvt_base6resultERNS_5rangeIKcLb1EEERNS3_IT_Lb1EEEmSt12codecvt_modeNS_10surrogatesE _ZNKSt7codecvtIDsciE5do_inERiPKcS3_RS3_PDsS5_RS5_ _ZNKSt25__codecvt_utf8_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ _ZNKSt19__codecvt_utf8_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ _ZNKSt19__codecvt_utf8_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ _ZNKSt19__codecvt_utf8_baseIDiE9do_lengthERiPKcS3_y _ZNSt12_GLOBAL__N_17ucs4_inERNS_5rangeIKcLb1EEERNS0_IDiLb1EEEmSt12codecvt_mode _ZNKSt7codecvtIDiciE5do_inERiPKcS3_RS3_PDiS5_RS5_ _ZNKSt19__codecvt_utf8_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ _ZNKSt20__codecvt_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ _ZNKSt7codecvtIDiciE9do_lengthERiPKcS3_y _ZNKSt7codecvtIDiciE6do_outERiPKDiS3_RS3_PcS5_RS5_ .rdata$_ZTSSt12co<      decvt_base .rdata$_ZTISt12codecvt_base .rdata$_ZTSSt23__codecvt_abstract_baseIwciE .rdata$_ZTISt23__codecvt_abstract_baseIwciE .rdata$_ZTSSt7codecvtIwciE .rdata$_ZTISt7codecvtIwciE .rdata$_ZTSSt23__codecvt_abstract_baseIDsciE .rdata$_ZTISt23__codecvt_abstract_baseIDsciE .rdata$_ZTSSt7codecvtIDsciE .rdata$_ZTISt7codecvtIDsciE .rdata$_ZTSSt23__codecvt_abstract_baseIDiciE .rdata$_ZTISt23__codecvt_abstract_baseIDiciE .rdata$_ZTSSt7codecvtIDiciE .rdata$_ZTISt7codecvtIDiciE .rdata$_ZTSSt19__codecvt_utf8_baseIDsE .rdata$_ZTISt19__codecvt_utf8_baseIDsE .rdata$_ZTSSt20__codecvt_utf16_baseIDsE .rdata$_ZTISt20__codecvt_utf16_baseIDsE .rdata$_ZTSSt25__codecvt_utf8_utf16_baseIDsE .rdata$_ZTISt25__codecvt_utf8_utf16_baseIDsE .rdata$_ZTSSt19__codecvt_utf8_baseIDiE .rdata$_ZTISt19__codecvt_utf8_baseIDiE .rdata$_ZTSSt20__codecvt_utf16_baseIDiE .rdata$_ZTISt20__codecvt_utf16_baseIDiE .rdata$_ZTSSt25__codecvt_utf8_utf16_baseIDiE .rdata$_ZTISt25__codecvt_utf8_utf16_baseIDiE .rdata$_ZTSSt19__codecvt_utf8_baseIwE .rdata$_Z=      TISt19__codecvt_utf8_baseIwE .rdata$_ZTSSt20__codecvt_utf16_baseIwE .rdata$_ZTISt20__codecvt_utf16_baseIwE .rdata$_ZTSSt25__codecvt_utf8_utf16_baseIwE .rdata$_ZTISt25__codecvt_utf8_utf16_baseIwE .rdata$_ZTVSt7codecvtIDsciE .rdata$_ZTVSt7codecvtIDiciE .rdata$_ZTVSt19__codecvt_utf8_baseIDsE .rdata$_ZTVSt19__codecvt_utf8_baseIDiE .rdata$_ZTVSt20__codecvt_utf16_baseIDsE .rdata$_ZTVSt20__codecvt_utf16_baseIDiE .rdata$_ZTVSt25__codecvt_utf8_utf16_baseIDsE .rdata$_ZTVSt25__codecvt_utf8_utf16_baseIDiE .text$_ZNSt12_GLOBAL__N_120read_utf8_code_pointERNS_5rangeIKcLb1EEEm .xdata$_ZNSt12_GLOBAL__N_120read_utf8_code_pointERNS_5rangeIKcLb1EEEm .pdata$_ZNSt12_GLOBAL__N_120read_utf8_code_pointERNS_5rangeIKcLb1EEEm .text$_ZNKSt7codecvtIDsciE10do_unshiftERiPcS2_RS2_ .xdata$_ZNKSt7codecvtIDsciE10do_unshiftERiPcS2_RS2_ .pdata$_ZNKSt7codecvtIDsciE10do_unshiftERiPcS2_RS2_ .text$_ZNKSt7codecvtIDsciE11do_encodingEv .xdata$_ZNKSt7codecvtIDsciE11do_encodingEv .pdata$_ZNKSt7codecvtIDsciE11do_encodingEv .text$_ZNKSt7codecvtIDsci>      E16do_always_noconvEv .xdata$_ZNKSt7codecvtIDsciE16do_always_noconvEv .pdata$_ZNKSt7codecvtIDsciE16do_always_noconvEv .text$_ZNKSt7codecvtIDsciE13do_max_lengthEv .xdata$_ZNKSt7codecvtIDsciE13do_max_lengthEv .pdata$_ZNKSt7codecvtIDsciE13do_max_lengthEv .text$_ZNKSt19__codecvt_utf8_baseIDsE13do_max_lengthEv .xdata$_ZNKSt19__codecvt_utf8_baseIDsE13do_max_lengthEv .pdata$_ZNKSt19__codecvt_utf8_baseIDsE13do_max_lengthEv .text$_ZNKSt19__codecvt_utf8_baseIDiE13do_max_lengthEv .xdata$_ZNKSt19__codecvt_utf8_baseIDiE13do_max_lengthEv .pdata$_ZNKSt19__codecvt_utf8_baseIDiE13do_max_lengthEv .text$_ZNKSt19__codecvt_utf8_baseIwE13do_max_lengthEv .xdata$_ZNKSt19__codecvt_utf8_baseIwE13do_max_lengthEv .pdata$_ZNKSt19__codecvt_utf8_baseIwE13do_max_lengthEv .text$_ZNKSt20__codecvt_utf16_baseIDsE13do_max_lengthEv .xdata$_ZNKSt20__codecvt_utf16_baseIDsE13do_max_lengthEv .pdata$_ZNKSt20__codecvt_utf16_baseIDsE13do_max_lengthEv .text$_ZNKSt20__codecvt_utf16_baseIDiE13do_max_lengthEv .xdata$_ZNKSt20__codecvt_utf16_baseIDiE1?      3do_max_lengthEv .pdata$_ZNKSt20__codecvt_utf16_baseIDiE13do_max_lengthEv .text$_ZNKSt20__codecvt_utf16_baseIwE13do_max_lengthEv .xdata$_ZNKSt20__codecvt_utf16_baseIwE13do_max_lengthEv .pdata$_ZNKSt20__codecvt_utf16_baseIwE13do_max_lengthEv .text$_ZNKSt25__codecvt_utf8_utf16_baseIDsE13do_max_lengthEv .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE13do_max_lengthEv .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE13do_max_lengthEv .text$_ZNKSt25__codecvt_utf8_utf16_baseIDiE13do_max_lengthEv .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE13do_max_lengthEv .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE13do_max_lengthEv .text$_ZNKSt25__codecvt_utf8_utf16_baseIwE13do_max_lengthEv .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE13do_max_lengthEv .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE13do_max_lengthEv .text$_ZNSt7codecvtIDsciED2Ev .xdata$_ZNSt7codecvtIDsciED2Ev .pdata$_ZNSt7codecvtIDsciED2Ev .text$_ZNSt19__codecvt_utf8_baseIDsED2Ev .xdata$_ZNSt19__codecvt_utf8_baseIDsED2Ev .pdata$_ZNSt19__codecvt_utf8_baseIDsED2Ev .text$@      _ZNSt20__codecvt_utf16_baseIDsED2Ev .xdata$_ZNSt20__codecvt_utf16_baseIDsED2Ev .pdata$_ZNSt20__codecvt_utf16_baseIDsED2Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIDsED2Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIDsED2Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIDsED2Ev .text$_ZNSt7codecvtIDiciED2Ev .xdata$_ZNSt7codecvtIDiciED2Ev .pdata$_ZNSt7codecvtIDiciED2Ev .text$_ZNSt19__codecvt_utf8_baseIDiED2Ev .xdata$_ZNSt19__codecvt_utf8_baseIDiED2Ev .pdata$_ZNSt19__codecvt_utf8_baseIDiED2Ev .text$_ZNSt20__codecvt_utf16_baseIDiED2Ev .xdata$_ZNSt20__codecvt_utf16_baseIDiED2Ev .pdata$_ZNSt20__codecvt_utf16_baseIDiED2Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIDiED2Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIDiED2Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIDiED2Ev .text$_ZNSt7codecvtIDsciED0Ev .xdata$_ZNSt7codecvtIDsciED0Ev .pdata$_ZNSt7codecvtIDsciED0Ev .text$_ZNSt19__codecvt_utf8_baseIDsED0Ev .xdata$_ZNSt19__codecvt_utf8_baseIDsED0Ev .pdata$_ZNSt19__codecvt_utf8_baseIDsED0Ev .text$_ZNSt20__codecvt_utf16_baseIDsED0Ev .xdaA      ta$_ZNSt20__codecvt_utf16_baseIDsED0Ev .pdata$_ZNSt20__codecvt_utf16_baseIDsED0Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIDsED0Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIDsED0Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIDsED0Ev .text$_ZNSt7codecvtIDiciED0Ev .xdata$_ZNSt7codecvtIDiciED0Ev .pdata$_ZNSt7codecvtIDiciED0Ev .text$_ZNSt19__codecvt_utf8_baseIDiED0Ev .xdata$_ZNSt19__codecvt_utf8_baseIDiED0Ev .pdata$_ZNSt19__codecvt_utf8_baseIDiED0Ev .text$_ZNSt20__codecvt_utf16_baseIDiED0Ev .xdata$_ZNSt20__codecvt_utf16_baseIDiED0Ev .pdata$_ZNSt20__codecvt_utf16_baseIDiED0Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIDiED0Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIDiED0Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIDiED0Ev .text$_ZNSt12_GLOBAL__N_18read_bomIKDsLb0ELy2EEEbRNS_5rangeIT_XT0_EEERAT1__Kh .xdata$_ZNSt12_GLOBAL__N_18read_bomIKDsLb0ELy2EEEbRNS_5rangeIT_XT0_EEERAT1__Kh .pdata$_ZNSt12_GLOBAL__N_18read_bomIKDsLb0ELy2EEEbRNS_5rangeIT_XT0_EEERAT1__Kh .text$_ZNSt12_GLOBAL__N_121read_utf16_code_pointILb0EEEDiRNS_5rangeB      IKDsXT_EEEmSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_121read_utf16_code_pointILb0EEEDiRNS_5rangeIKDsXT_EEEmSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_121read_utf16_code_pointILb0EEEDiRNS_5rangeIKDsXT_EEEmSt12codecvt_mode .text$_ZNSt19__codecvt_utf8_baseIwED2Ev .xdata$_ZNSt19__codecvt_utf8_baseIwED2Ev .pdata$_ZNSt19__codecvt_utf8_baseIwED2Ev .text$_ZNSt19__codecvt_utf8_baseIwED0Ev .xdata$_ZNSt19__codecvt_utf8_baseIwED0Ev .pdata$_ZNSt19__codecvt_utf8_baseIwED0Ev .text$_ZNSt20__codecvt_utf16_baseIwED2Ev .xdata$_ZNSt20__codecvt_utf16_baseIwED2Ev .pdata$_ZNSt20__codecvt_utf16_baseIwED2Ev .text$_ZNSt20__codecvt_utf16_baseIwED0Ev .xdata$_ZNSt20__codecvt_utf16_baseIwED0Ev .pdata$_ZNSt20__codecvt_utf16_baseIwED0Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIwED2Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIwED2Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIwED2Ev .text$_ZNSt25__codecvt_utf8_utf16_baseIwED0Ev .xdata$_ZNSt25__codecvt_utf8_utf16_baseIwED0Ev .pdata$_ZNSt25__codecvt_utf8_utf16_baseIwED0Ev .text$_ZNSt12_GLOBAL__C      N_121write_utf8_code_pointERNS_5rangeIcLb1EEEDi .xdata$_ZNSt12_GLOBAL__N_121write_utf8_code_pointERNS_5rangeIcLb1EEEDi .pdata$_ZNSt12_GLOBAL__N_121write_utf8_code_pointERNS_5rangeIcLb1EEEDi .text$_ZNSt12_GLOBAL__N_115write_utf16_bomILb0EEEbRNS_5rangeIDsXT_EEESt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_115write_utf16_bomILb0EEEbRNS_5rangeIDsXT_EEESt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_115write_utf16_bomILb0EEEbRNS_5rangeIDsXT_EEESt12codecvt_mode .text$_ZNKSt20__codecvt_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .pdata$_ZNKSt20__codecvt_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .text$_ZNSt12_GLOBAL__N_114write_utf8_bomERNS_5rangeIcLb1EEESt12codecvt_mode.part.19 .xdata$_ZNSt12_GLOBAL__N_114write_utf8_bomERNS_5rangeIcLb1EEESt12codecvt_mode.part.19 .pdata$_ZNSt12_GLOBAL__N_114write_utf8_bomERNS_5rangeIcLb1EEESt12codecvt_mode.part.19 .text$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSD      t12codecvt_modeNS_10surrogatesE.part.20 .xdata$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE.part.20 .pdata$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE.part.20 .text$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE .xdata$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE .pdata$_ZNSt12_GLOBAL__N_19utf16_outIDsEENSt12codecvt_base6resultERNS_5rangeIKT_Lb1EEERNS3_IcLb1EEEmSt12codecvt_modeNS_10surrogatesE .text$_ZNKSt25__codecvt_utf8_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .xdaE      ta$_ZNKSt19__codecvt_utf8_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .xdata$_ZNKSt19__codecvt_utf8_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .text$_ZNKSt7codecvtIDsciE6do_outERiPKDsS3_RS3_PcS5_RS5_ .xdata$_ZNKSt7codecvtIDsciE6do_outERiPKDsS3_RS3_PcS5_RS5_ .pdata$_ZNKSt7codecvtIDsciE6do_outERiPKDsS3_RS3_PcS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .xdata$_ZNKSt19__codecvt_utf8_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .text$_ZNSt12_GLOBAL__N_114read_utf16_bomILb0EEEvRNS_5rangeIKDsXT_EEERSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_114read_utf16_bomILb0EEEvRNS_5rangeIKDsXT_EEERSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_114read_utf16_bomILb0EEEvRNS_5rangeIKDsXT_EEERSt12codecvt_mode .text$_ZNKSt20__codecvt_utf16_baseIDiE5dF      o_inERiPKcS3_RS3_PDiS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .pdata$_ZNKSt20__codecvt_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .text$_ZNKSt20__codecvt_utf16_baseIDiE9do_lengthERiPKcS3_y .xdata$_ZNKSt20__codecvt_utf16_baseIDiE9do_lengthERiPKcS3_y .pdata$_ZNKSt20__codecvt_utf16_baseIDiE9do_lengthERiPKcS3_y .text$_ZNSt12_GLOBAL__N_17ucs2_inERNS_5rangeIKDsLb0EEERNS0_IDsLb1EEEDiSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_17ucs2_inERNS_5rangeIKDsLb0EEERNS0_IDsLb1EEEDiSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_17ucs2_inERNS_5rangeIKDsLb0EEERNS0_IDsLb1EEEDiSt12codecvt_mode .text$_ZNKSt20__codecvt_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .pdata$_ZNKSt20__codecvt_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .text$_ZNKSt20__codecvt_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .pdata$_ZNKSt20__codecvt_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .tG      ext$_ZNSt12_GLOBAL__N_19ucs2_spanERNS_5rangeIKDsLb0EEEyDiSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_19ucs2_spanERNS_5rangeIKDsLb0EEEyDiSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_19ucs2_spanERNS_5rangeIKDsLb0EEEyDiSt12codecvt_mode .text$_ZNKSt20__codecvt_utf16_baseIDsE9do_lengthERiPKcS3_y .xdata$_ZNKSt20__codecvt_utf16_baseIDsE9do_lengthERiPKcS3_y .pdata$_ZNKSt20__codecvt_utf16_baseIDsE9do_lengthERiPKcS3_y .text$_ZNKSt20__codecvt_utf16_baseIwE9do_lengthERiPKcS3_y .xdata$_ZNKSt20__codecvt_utf16_baseIwE9do_lengthERiPKcS3_y .pdata$_ZNKSt20__codecvt_utf16_baseIwE9do_lengthERiPKcS3_y .text$_ZNSt12_GLOBAL__N_18ucs2_outERNS_5rangeIKDsLb1EEERNS0_IDsLb0EEEDiSt12codecvt_mode.part.23 .xdata$_ZNSt12_GLOBAL__N_18ucs2_outERNS_5rangeIKDsLb1EEERNS0_IDsLb0EEEDiSt12codecvt_mode.part.23 .pdata$_ZNSt12_GLOBAL__N_18ucs2_outERNS_5rangeIKDsLb1EEERNS0_IDsLb0EEEDiSt12codecvt_mode.part.23 .text$_ZNKSt20__codecvt_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .pdaH      ta$_ZNKSt20__codecvt_utf16_baseIDsE6do_outERiPKDsS3_RS3_PcS5_RS5_ .text$_ZNKSt25__codecvt_utf8_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .text$_ZNKSt25__codecvt_utf8_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE6do_outERiPKDiS3_RS3_PcS5_RS5_ .text$_ZNSt12_GLOBAL__N_18read_bomIKcLb1ELy3EEEbRNS_5rangeIT_XT0_EEERAT1__Kh.constprop.29 .xdata$_ZNSt12_GLOBAL__N_18read_bomIKcLb1ELy3EEEbRNS_5rangeIT_XT0_EEERAT1__Kh.constprop.29 .pdata$_ZNSt12_GLOBAL__N_18read_bomIKcLb1ELy3EEEbRNS_5rangeIT_XT0_EEERAT1__Kh.constprop.29 .text$_ZNKSt25__codecvt_utf8_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .text$_ZNKSt25_I      _codecvt_utf8_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .text$_ZNSt12_GLOBAL__N_19ucs2_spanEPKcS1_yDiSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_19ucs2_spanEPKcS1_yDiSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_19ucs2_spanEPKcS1_yDiSt12codecvt_mode .text$_ZNKSt19__codecvt_utf8_baseIDsE9do_lengthERiPKcS3_y .xdata$_ZNKSt19__codecvt_utf8_baseIDsE9do_lengthERiPKcS3_y .pdata$_ZNKSt19__codecvt_utf8_baseIDsE9do_lengthERiPKcS3_y .text$_ZNKSt19__codecvt_utf8_baseIwE9do_lengthERiPKcS3_y .xdata$_ZNKSt19__codecvt_utf8_baseIwE9do_lengthERiPKcS3_y .pdata$_ZNKSt19__codecvt_utf8_baseIwE9do_lengthERiPKcS3_y .text$_ZNSt12_GLOBAL__N_110utf16_spanEPKcS1_yDiSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_110utf16_spanEPKcS1_yDiSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_110utf16_spanEPKcS1_yDiSt12codecvt_mode .text$_ZNKSt7codecvtIDsciE9do_lengthERiPKcS3_y .xdata$_ZNKSt7codecvtIDsciE9do_lengthEJ      RiPKcS3_y .pdata$_ZNKSt7codecvtIDsciE9do_lengthERiPKcS3_y .text$_ZNKSt25__codecvt_utf8_utf16_baseIDsE9do_lengthERiPKcS3_y .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE9do_lengthERiPKcS3_y .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE9do_lengthERiPKcS3_y .text$_ZNKSt25__codecvt_utf8_utf16_baseIDiE9do_lengthERiPKcS3_y .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE9do_lengthERiPKcS3_y .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDiE9do_lengthERiPKcS3_y .text$_ZNKSt25__codecvt_utf8_utf16_baseIwE9do_lengthERiPKcS3_y .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE9do_lengthERiPKcS3_y .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIwE9do_lengthERiPKcS3_y .text$_ZNSt12_GLOBAL__N_18utf16_inIDsEENSt12codecvt_base6resultERNS_5rangeIKcLb1EEERNS3_IT_Lb1EEEmSt12codecvt_modeNS_10surrogatesE .xdata$_ZNSt12_GLOBAL__N_18utf16_inIDsEENSt12codecvt_base6resultERNS_5rangeIKcLb1EEERNS3_IT_Lb1EEEmSt12codecvt_modeNS_10surrogatesE .pdata$_ZNSt12_GLOBAL__N_18utf16_inIDsEENSt12codecvt_base6resultERNS_5rangeIKcLb1EEERNS3_IT_Lb1EEEmSt12codecvt_modeNK      S_10surrogatesE .text$_ZNKSt7codecvtIDsciE5do_inERiPKcS3_RS3_PDsS5_RS5_ .xdata$_ZNKSt7codecvtIDsciE5do_inERiPKcS3_RS3_PDsS5_RS5_ .pdata$_ZNKSt7codecvtIDsciE5do_inERiPKcS3_RS3_PDsS5_RS5_ .text$_ZNKSt25__codecvt_utf8_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .xdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .pdata$_ZNKSt25__codecvt_utf8_utf16_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .xdata$_ZNKSt19__codecvt_utf8_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIDsE5do_inERiPKcS3_RS3_PDsS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .xdata$_ZNKSt19__codecvt_utf8_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIwE5do_inERiPKcS3_RS3_PwS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIDiE9do_lengthERiPKcS3_y .xdata$_ZNKSt19__codecvt_utf8_baseIDiE9do_lengthERiPKcS3_y .pdata$_ZNKSt19__codecvt_utf8_baseIDiE9do_lengthERiPKcS3_y .text$_ZNSt12_GLOBAL__N_17ucs4_inL      ERNS_5rangeIKcLb1EEERNS0_IDiLb1EEEmSt12codecvt_mode .xdata$_ZNSt12_GLOBAL__N_17ucs4_inERNS_5rangeIKcLb1EEERNS0_IDiLb1EEEmSt12codecvt_mode .pdata$_ZNSt12_GLOBAL__N_17ucs4_inERNS_5rangeIKcLb1EEERNS0_IDiLb1EEEmSt12codecvt_mode .text$_ZNKSt7codecvtIDiciE5do_inERiPKcS3_RS3_PDiS5_RS5_ .xdata$_ZNKSt7codecvtIDiciE5do_inERiPKcS3_RS3_PDiS5_RS5_ .pdata$_ZNKSt7codecvtIDiciE5do_inERiPKcS3_RS3_PDiS5_RS5_ .text$_ZNKSt19__codecvt_utf8_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .xdata$_ZNKSt19__codecvt_utf8_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .pdata$_ZNKSt19__codecvt_utf8_baseIDiE5do_inERiPKcS3_RS3_PDiS5_RS5_ .text$_ZNKSt20__codecvt_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .xdata$_ZNKSt20__codecvt_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .pdata$_ZNKSt20__codecvt_utf16_baseIwE6do_outERiPKwS3_RS3_PcS5_RS5_ .text$_ZNKSt7codecvtIDiciE9do_lengthERiPKcS3_y .xdata$_ZNKSt7codecvtIDiciE9do_lengthERiPKcS3_y .pdata$_ZNKSt7codecvtIDiciE9do_lengthERiPKcS3_y .text$_ZNKSt7codecvtIDiciE6do_outERiPKDiS3_RS3_PcS5_RS5_ .xdata$_ZNKSt7coM      decvtIDiciE6do_outERiPKDiS3_RS3_PcS5_RS5_ .pdata$_ZNKSt7codecvtIDiciE6do_outERiPKDiS3_RS3_PcS5_RS5_ .data$_ZNSt7codecvtIDiciE2idE .data$_ZNSt7codecvtIDsciE2idE .rdata$_ZNSt12_GLOBAL__N_1L11utf16le_bomE .rdata$_ZNSt12_GLOBAL__N_1L9utf16_bomE .rdata$_ZNSt12_GLOBAL__N_1L8utf8_bomE _ZNSt6locale5_Impl13_M_init_extraEPPNS_5facetE _ZNSt12_GLOBAL__N_110numpunct_cE .rdata$.refptr._ZNSt8numpunctIcE2idE .rdata$.refptr._ZTVSt7collateIcE _ZNSt12_GLOBAL__N_19collate_cE .rdata$.refptr._ZNSt7collateIcE2idE _ZNSt12_GLOBAL__N_113moneypunct_cfE .rdata$.refptr._ZNSt10moneypunctIcLb0EE2idE _ZNSt12_GLOBAL__N_113moneypunct_ctE .rdata$.refptr._ZNSt10moneypunctIcLb1EE2idE .rdata$.refptr._ZTVSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt12_GLOBAL__N_111money_get_cE .rdata$.refptr._ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt12_GLOBAL__N_111money_put_cE .rdata$.refptr._ZNSt9money_putIcSt19ostreambuf_iteraN      torIcSt11char_traitsIcEEE2idE .rdata$.refptr._ZTVSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt12_GLOBAL__N_110time_get_cE .rdata$.refptr._ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt12_GLOBAL__N_110messages_cE .rdata$.refptr._ZNSt8messagesIcE2idE _ZNSt12_GLOBAL__N_110numpunct_wE .rdata$.refptr._ZNSt8numpunctIwE2idE .rdata$.refptr._ZTVSt7collateIwE _ZNSt12_GLOBAL__N_19collate_wE .rdata$.refptr._ZNSt7collateIwE2idE _ZNSt12_GLOBAL__N_113moneypunct_wfE .rdata$.refptr._ZNSt10moneypunctIwLb0EE2idE _ZNSt12_GLOBAL__N_113moneypunct_wtE .rdata$.refptr._ZNSt10moneypunctIwLb1EE2idE .rdata$.refptr._ZTVSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt12_GLOBAL__N_111money_get_wE .rdata$.refptr._ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$.refptr._ZTVSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt12_GLOBAL__N_111money_put_wE .rdata$.refptr._ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdaO      ta$.refptr._ZTVSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt12_GLOBAL__N_110time_get_wE .rdata$.refptr._ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZNSt12_GLOBAL__N_110messages_wE .rdata$.refptr._ZNSt8messagesIwE2idE _ZNSt6locale5_Impl13_M_init_extraEPvS1_PKcS3_ _ZNKSt6locale4nameEv .text$_ZNSt6locale5_Impl13_M_init_extraEPPNS_5facetE .xdata$_ZNSt6locale5_Impl13_M_init_extraEPPNS_5facetE .pdata$_ZNSt6locale5_Impl13_M_init_extraEPPNS_5facetE .text$_ZNSt6locale5_Impl13_M_init_extraEPvS1_PKcS3_ .xdata$_ZNSt6locale5_Impl13_M_init_extraEPvS1_PKcS3_ .pdata$_ZNSt6locale5_Impl13_M_init_extraEPvS1_PKcS3_ .text$_ZNKSt6locale4nameEv .xdata$_ZNKSt6locale4nameEv .pdata$_ZNKSt6locale4nameEv .data$_ZNSt12_GLOBAL__N_110messages_wE .data$_ZNSt12_GLOBAL__N_110time_get_wE .data$_ZNSt12_GLOBAL__N_111money_put_wE .data$_ZNSt12_GLOBAL__N_111money_get_wE .data$_ZNSt12_GLOBAL__N_113moneypunct_wfE .data$_ZNSt12_GLOBAL__N_113moneypunct_wtE .data$_ZNSt12_GLOBAL__N_110numpunct_wE .data$_ZP      NSt12_GLOBAL__N_19collate_wE .data$_ZNSt12_GLOBAL__N_110messages_cE .data$_ZNSt12_GLOBAL__N_110time_get_cE .data$_ZNSt12_GLOBAL__N_111money_put_cE .data$_ZNSt12_GLOBAL__N_111money_get_cE .data$_ZNSt12_GLOBAL__N_113moneypunct_cfE .data$_ZNSt12_GLOBAL__N_113moneypunct_ctE .data$_ZNSt12_GLOBAL__N_110numpunct_cE .data$_ZNSt12_GLOBAL__N_19collate_cE _ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE10do_compareEPKcS4_S4_S4_ _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_yearESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE16do_get_monthnameESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE14do_get_weekdayESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_dateESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IosQ      tateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_timeESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE13do_date_orderEv _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basece _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE8do_closeEi _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKSsRKSt6locale _ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE10do_compareEPKwS4_S4_S4_ _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_yearESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE16do_get_monthnameESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZR      NKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE14do_get_weekdayESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_dateESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_timeESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE13do_date_orderEv _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewe _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE8do_closeEi _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKSsRKSt6locale _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11chS      ar_traitsIwEEbRSt8ios_basewRKSbIwS5_SaIwEE _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKSs _ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE12do_transformEPKwS4_ _ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE12do_transformEPKcS4_ _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKSs _ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIwEEvPv _ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIcEEvPv _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED2Ev _ZTVNSt13__facet_shT      ims12_GLOBAL__N_113time_get_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED2Ev _ZTU      VNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED1Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED1Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED1Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_V      shimIwLb1EED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED0Ev _ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED1Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED0Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED2Ev _ZTVNSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED1Ev _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED0Ev _ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED0Ev _ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED0Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED0Ev _ZNSt13__facet_shims12_GLOBALW      __N_115moneypunct_shimIwLb1EED0Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED0Ev _ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED0Ev _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED0Ev _ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED0Ev _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRSbIwS5_SaIwEE _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt6locale5facet19_M_remove_referenceEv _ZNKSt6locale5facet19_M_remove_referenceEv .text$_ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E _ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .text$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16_X      _numpunct_cacheIT_E _ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .text$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ _ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .text$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ _ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .text$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ _ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .text$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ _ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLbY      0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNStZ      13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ _ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .text$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ _ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .text$_ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y _ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .text$_ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y _ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .te[      xt$_ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi _ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .text$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi _ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .text$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE _ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .text$_ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE _ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .text$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseR\      St12_Ios_IostateP2tmc _ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .text$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc _ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .text$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE _ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EES]      t17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE _ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE _ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE _ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE _ZNKSt6locale5facet11_M^      _cow_shimEPKNS_2idE .rdata$_ZTINSt6locale5facet6__shimE _ZTINSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE _ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE _ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE _ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE _ZTINSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE _ZTINSt13__facet_shims12_GLOBAL__N_112_      collate_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE _ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE _ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE _ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE _ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE _ZTINSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE _ZTINSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE _ZTINSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE .rdata$_ZTSNSt6locale5facet6__shimE _ZTINSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE _ZTSNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE _ZTINSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE _ZTSNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE10do_compareEPKcS4_S4_S4_ .xdata$_ZNKS`      t13__facet_shims12_GLOBAL__N_112collate_shimIcE10do_compareEPKcS4_S4_S4_ .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE10do_compareEPKcS4_S4_S4_ .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_yearESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_yearESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_yearESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE16do_get_monthnameESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE16do_get_monthnameESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE16do_get_monthna      ameESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE14do_get_weekdayESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE14do_get_weekdayESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE14do_get_weekdayESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_dateESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_dateESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_dateESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_Iostatb      eP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_timeESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_timeESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE11do_get_timeESt19istreambuf_iteratorIcSt11char_traitsIcEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE13do_date_orderEv .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE13do_date_orderEv .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIcE13do_date_orderEv .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt13_c      _facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basece .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basece .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basece .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE8do_closeEi .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE8do_closeEi .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE8do_closeEi .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKSsRKSt6locale .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKSsRKSt6locale .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKSsRKSt6locale .text$_ZNKSt13__facet_shims1d      2_GLOBAL__N_112collate_shimIwE10do_compareEPKwS4_S4_S4_ .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE10do_compareEPKwS4_S4_S4_ .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE10do_compareEPKwS4_S4_S4_ .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_yearESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_yearESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_yearESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE16do_get_monthnameESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE16do_get_monthnameESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$e      _ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE16do_get_monthnameESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE14do_get_weekdayESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE14do_get_weekdayESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE14do_get_weekdayESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_dateESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_dateESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_dateESt19istf      reambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_timeESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_timeESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE11do_get_timeESt19istreambuf_iteratorIwSt11char_traitsIwEES6_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE13do_date_orderEv .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE13do_date_orderEv .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113time_get_shimIwE13do_date_orderEv .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt1g      1char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewe .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewe .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewe .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE8do_closeEi .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE8do_closeEi .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE8do_closeEi .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKSsRKSt6locale .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKSsRKSt6locale .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113mh      essages_shimIwE7do_openERKSsRKSt6locale .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKSbIwS5_SaIwEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKSbIwS5_SaIwEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKSbIwS5_SaIwEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKSs .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKSs .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKSs .text$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE12do_transformEPKwS4_ .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE12do_transformi      EPKwS4_ .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIwE12do_transformEPKwS4_ .text$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE12do_transformEPKcS4_ .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE12do_transformEPKcS4_ .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_112collate_shimIcE12do_transformEPKcS4_ .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKSs .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKSs .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKSs .text$_ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIwEEvPv .xdata$_ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIwEEvPv .pdata$_ZNSt13__facej      t_shims12_GLOBAL__N_116__destroy_stringIwEEvPv .text$_ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIcEEvPv .xdata$_ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIcEEvPv .pdata$_ZNSt13__facet_shims12_GLOBAL__N_116__destroy_stringIcEEvPv .text$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED2Ev .textk      $_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shil      mIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113tm      ime_get_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL_n      _N_114money_get_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED2Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED2Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED2Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIwED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113messages_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLo      OBAL__N_113numpunct_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EED0Ev .pdata$_ZNSt13__facet_shimsp      12_GLOBAL__N_115moneypunct_shimIwLb0EED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIcED0Ev .text$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED0Ev .xdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED0Ev .pdata$_ZNSt13__facet_shims12_GLOBAL__N_112collate_shimIwED0Ev .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRSbIwS5_SaIwEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRSbIwS5_SaIwEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRSbIwS5_SaIwEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_q      bRSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt6locale5facet19_M_remove_referenceEv .pdata$_ZNKSt6locale5facet19_M_remove_referenceEv .xdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .pdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .xdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .pdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .xdata$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constar      ntIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .pdata$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .xdata$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .pdata$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKT_S9_S9_S9_ .xdata$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .pdata$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .xdata$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .pdata$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cachs      eIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__fat      cet_shims15__messages_openIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .pdata$_ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .xdata$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .pdata$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb0EEPKNSt6locale5facetEPKcyRKS3_ .xdata$_ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .pdata$_ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .xdata$_ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .pdata$_ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .xdata$_ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .pdata$_ZNSt13__facu      et_shims16__messages_closeIcEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .xdata$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .pdata$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb0EEPKNSt6locale5facetEi .xdata$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .pdata$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .xdata$_ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .pdata$_ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb0EEPKNSt6locale5facetE .xdata$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .pdata$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_itv      eratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .xdata$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .pdata$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .xdata$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8iw      os_baseRSt12_Ios_IostatePePNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb0EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .text$_ZNKSt6locale5facet11_M_cow_shimEPKNS_2idE .xdata$_Zx      NKSt6locale5facet11_M_cow_shimEPKNS_2idE .pdata$_ZNKSt6locale5facet11_M_cow_shimEPKNS_2idE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE .rdata$_ZTINSt13_y      _facet_shims12_GLOBAL__N_113numpunct_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113messages_shimIwEE .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEEz       .rdata$_ZTINSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE .rdata$_ZTSNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_112collate_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb1EEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIcLb0EEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_114money_get_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_114money_put_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_113messages_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_113numpunct_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_112collate_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb1EEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_115moneypunct_shimIwLb0EEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_114money_get_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_114money_put_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_11{      3messages_shimIwEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_113time_get_shimIcEE .rdata$_ZTVNSt13__facet_shims12_GLOBAL__N_113time_get_shimIwEE .text$_ZNKSs7_M_dataEv _ZNKSs7_M_dataEv .text$_ZNSs7_M_dataEPc _ZNSs7_M_dataEPc .text$_ZNKSs6_M_repEv _ZNKSs6_M_repEv .text$_ZNKSs9_M_ibeginEv _ZNKSs9_M_ibeginEv .text$_ZNKSs7_M_iendEv _ZNKSs7_M_iendEv .text$_ZNKSs8_M_checkEyPKc _ZNKSs8_M_checkEyPKc .text$_ZNKSs15_M_check_lengthEyyPKc _ZNKSs15_M_check_lengthEyyPKc .text$_ZNKSs8_M_limitEyy _ZNKSs8_M_limitEyy .text$_ZNKSs11_M_disjunctEPKc _ZNKSs11_M_disjunctEPKc .text$_ZNSs7_M_copyEPcPKcy _ZNSs7_M_copyEPcPKcy .text$_ZNSs7_M_moveEPcPKcy _ZNSs7_M_moveEPcPKcy .text$_ZNSs9_M_assignEPcyc _ZNSs9_M_assignEPcyc .text$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ .text$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ .text$_ZNSs13_S_copy_charsEPcS_S_ _ZNSs13_S|      _copy_charsEPcS_S_ .text$_ZNSs13_S_copy_charsEPcPKcS1_ _ZNSs13_S_copy_charsEPcPKcS1_ .text$_ZNSs10_S_compareEyy _ZNSs10_S_compareEyy .text$_ZNSs12_S_empty_repEv _ZNSs12_S_empty_repEv .data$_ZNSs4_Rep20_S_empty_rep_storageE .text$_ZNSsD2Ev _ZNSsD2Ev .text$_ZNSsD1Ev _ZNSsD1Ev .text$_ZNKSs5beginEv _ZNKSs5beginEv .text$_ZNKSs3endEv _ZNKSs3endEv .text$_ZNKSs6rbeginEv _ZNKSs6rbeginEv .text$_ZNKSs4rendEv _ZNKSs4rendEv .text$_ZNKSs6cbeginEv _ZNKSs6cbeginEv .text$_ZNKSs4cendEv _ZNKSs4cendEv .text$_ZNKSs7crbeginEv _ZNKSs7crbeginEv .text$_ZNKSs5crendEv _ZNKSs5crendEv .text$_ZNKSs4sizeEv _ZNKSs4sizeEv .text$_ZNKSs6lengthEv _ZNKSs6lengthEv .text$_ZNKSs8max_sizeEv _ZNKSs8max_sizeEv .text$_ZNKSs8capacityEv _ZNKSs8capacityEv .text$_ZNKSs5emptyEv _ZNKSs5emptyEv .text$_ZNKSsixEy _ZNKSsixEy .text$_ZNKSs2atEy _ZNKSs2atEy .text$_ZNKSs5frontEv _ZNKSs5frontEv .text$_ZNKSs4backEv _ZNKSs4backEv .text$_ZNKSs4copyEPcyy _ZNKSs4copyEPcyy .text$_ZNSs4swapERSs _ZNSs4swapERSs .text$_ZNSsaSEOSs _ZNSsaSEOSs .text$_ZNSs6assignEOSs _ZNS}      s6assignEOSs .text$_ZNKSs5c_strEv _ZNKSs5c_strEv .text$_ZNKSs4dataEv _ZNKSs4dataEv .text$_ZNKSs13get_allocatorEv _ZNKSs13get_allocatorEv .text$_ZNKSs4findEPKcyy _ZNKSs4findEPKcyy .text$_ZNKSs4findERKSsy _ZNKSs4findERKSsy .text$_ZNKSs4findEPKcy _ZNKSs4findEPKcy .text$_ZNKSs4findEcy _ZNKSs4findEcy .text$_ZNKSs5rfindEPKcyy _ZNKSs5rfindEPKcyy .text$_ZNKSs5rfindERKSsy _ZNKSs5rfindERKSsy .text$_ZNKSs5rfindEPKcy _ZNKSs5rfindEPKcy .text$_ZNKSs5rfindEcy _ZNKSs5rfindEcy .text$_ZNKSs13find_first_ofEPKcyy _ZNKSs13find_first_ofEPKcyy .text$_ZNKSs13find_first_ofERKSsy _ZNKSs13find_first_ofERKSsy .text$_ZNKSs13find_first_ofEPKcy _ZNKSs13find_first_ofEPKcy .text$_ZNKSs13find_first_ofEcy _ZNKSs13find_first_ofEcy .text$_ZNKSs12find_last_ofEPKcyy _ZNKSs12find_last_ofEPKcyy .text$_ZNKSs12find_last_ofERKSsy _ZNKSs12find_last_ofERKSsy .text$_ZNKSs12find_last_ofEPKcy _ZNKSs12find_last_ofEPKcy .text$_ZNKSs12find_last_ofEcy _ZNKSs12find_last_ofEcy .text$_ZNKSs17find_first_not_ofEPKcyy _ZNKSs17find_first_not_ofEPKcyy .text$_ZN~      KSs17find_first_not_ofERKSsy _ZNKSs17find_first_not_ofERKSsy .text$_ZNKSs17find_first_not_ofEPKcy _ZNKSs17find_first_not_ofEPKcy .text$_ZNKSs17find_first_not_ofEcy _ZNKSs17find_first_not_ofEcy .text$_ZNKSs16find_last_not_ofEPKcyy _ZNKSs16find_last_not_ofEPKcyy .text$_ZNKSs16find_last_not_ofERKSsy _ZNKSs16find_last_not_ofERKSsy .text$_ZNKSs16find_last_not_ofEPKcy _ZNKSs16find_last_not_ofEPKcy .text$_ZNKSs16find_last_not_ofEcy _ZNKSs16find_last_not_ofEcy .text$_ZNKSs7compareERKSs _ZNKSs7compareERKSs .text$_ZNKSs7compareEyyRKSs _ZNKSs7compareEyyRKSs .text$_ZNKSs7compareEyyRKSsyy _ZNKSs7compareEyyRKSsyy .text$_ZNKSs7compareEPKc _ZNKSs7compareEPKc .text$_ZNKSs7compareEyyPKc _ZNKSs7compareEyyPKc .text$_ZNKSs7compareEyyPKcy _ZNKSs7compareEyyPKcy .text$_ZNSs12_Alloc_hiderC2EPcRKSaIcE _ZNSs12_Alloc_hiderC2EPcRKSaIcE .text$_ZNSs12_Alloc_hiderC1EPcRKSaIcE _ZNSs12_Alloc_hiderC1EPcRKSaIcE .text$_ZNSs4_Rep12_S_empty_repEv _ZNSs4_Rep12_S_empty_repEv .text$_ZNKSs4_Rep12_M_is_leakedEv _ZNKSs4_Rep12_M_is_leakedEv .text      $_ZNKSs4_Rep12_M_is_sharedEv _ZNKSs4_Rep12_M_is_sharedEv .text$_ZNSs4_Rep13_M_set_leakedEv _ZNSs4_Rep13_M_set_leakedEv .text$_ZNSs4_Rep15_M_set_sharableEv _ZNSs4_Rep15_M_set_sharableEv .text$_ZNSs4_Rep26_M_set_length_and_sharableEy _ZNSs4_Rep26_M_set_length_and_sharableEy .text$_ZNSs4_Rep10_M_refdataEv _ZNSs4_Rep10_M_refdataEv .text$_ZNSs4_Rep9_S_createEyyRKSaIcE _ZNSs4_Rep9_S_createEyyRKSaIcE .text$_ZNSs9_M_mutateEyyy _ZNSs9_M_mutateEyyy .text$_ZNSs12_M_leak_hardEv _ZNSs12_M_leak_hardEv .text$_ZNSs7_M_leakEv _ZNSs7_M_leakEv .text$_ZNSs4rendEv _ZNSs4rendEv .text$_ZNSs5frontEv _ZNSs5frontEv .text$_ZNSsixEy _ZNSsixEy .text$_ZNSs5beginEv _ZNSs5beginEv .text$_ZNSs6rbeginEv _ZNSs6rbeginEv .text$_ZNSs3endEv _ZNSs3endEv .text$_ZNSs4backEv _ZNSs4backEv .text$_ZNSs2atEy _ZNSs2atEy .text$_ZNSs5clearEv _ZNSs5clearEv .text$_ZNSs5eraseEyy _ZNSs5eraseEyy .text$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE .text$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEES2�      _ _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEES2_ .text$_ZNSs14_M_replace_auxEyyyc _ZNSs14_M_replace_auxEyyyc .text$_ZNSs6assignEyc _ZNSs6assignEyc .text$_ZNSsaSEc _ZNSsaSEc .text$_ZNSs6insertEyyc _ZNSs6insertEyyc .text$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc .text$_ZNSs7replaceEyyyc _ZNSs7replaceEyyyc .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_yc _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_yc .text$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEyc _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEyc .text$_ZNSs15_M_replace_safeEyyPKcy _ZNSs15_M_replace_safeEyyPKcy .text$_ZNSs6assignEPKcy _ZNSs6assignEPKcy .text$_ZNSsaSESt16initializer_listIcE _ZNSsaSESt16initializer_listIcE .text$_ZNSs6assignERKSsyy _ZNSs6assignERKSsyy .text$_ZNSs6assignEPKc _ZNSs6assignEPKc .text$_ZNSsaSEPKc _ZNSsaSEPKc .text$_ZNSs6assignESt16initializer_listIcE _ZNSs6assignESt16initializer_listIcE .text$_ZNSs6insertEyPKcy _ZNSs6insert�      EyPKcy .text$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE .text$_ZNSs6insertEyRKSsyy _ZNSs6insertEyRKSsyy .text$_ZNSs6insertEyPKc _ZNSs6insertEyPKc .text$_ZNSs6insertEyRKSs _ZNSs6insertEyRKSs .text$_ZNSs8pop_backEv _ZNSs8pop_backEv .text$_ZNSs12_S_constructEycRKSaIcE _ZNSs12_S_constructEycRKSaIcE .text$_ZNSsC2Ev _ZNSsC2Ev .text$_ZNSsC1Ev _ZNSsC1Ev .text$_ZNSsC2ERKSaIcE _ZNSsC2ERKSaIcE .text$_ZNSsC1ERKSaIcE _ZNSsC1ERKSaIcE .text$_ZNSsC2EycRKSaIcE _ZNSsC2EycRKSaIcE .text$_ZNSsC1EycRKSaIcE _ZNSsC1EycRKSaIcE .text$_ZNSsC2EOSs _ZNSsC2EOSs .text$_ZNSsC1EOSs _ZNSsC1EOSs .text$_ZNSs18_S_construct_aux_2EycRKSaIcE _ZNSs18_S_construct_aux_2EycRKSaIcE .text$_ZNSs4_Rep10_M_disposeERKSaIcE _ZNSs4_Rep10_M_disposeERKSaIcE .text$_ZNSs4_Rep10_M_destroyERKSaIcE _ZNSs4_Rep10_M_destroyERKSaIcE .text$_ZNSs4_Rep10_M_refcopyEv _ZNSs4_Rep10_M_refcopyEv .text$_ZNSs4_Rep8_M_cloneERKSaIcEy _ZNSs4_Rep8_M_cloneERKSaIcEy .text$_ZN�      Ss7reserveEy _ZNSs7reserveEy .text$_ZNSs13shrink_to_fitEv _ZNSs13shrink_to_fitEv .text$_ZNSs6appendERKSs _ZNSs6appendERKSs .text$_ZNSspLERKSs _ZNSspLERKSs .text$_ZNSs6appendERKSsyy _ZNSs6appendERKSsyy .text$_ZNSs6appendEPKcy _ZNSs6appendEPKcy .text$_ZNSspLESt16initializer_listIcE _ZNSspLESt16initializer_listIcE .text$_ZNSs6appendEPKc _ZNSs6appendEPKc .text$_ZNSspLEPKc _ZNSspLEPKc .text$_ZNSs6appendESt16initializer_listIcE _ZNSs6appendESt16initializer_listIcE _ZNSs6appendEyc.part.20 .text$_ZNSs6appendEyc _ZNSs6appendEyc .text$_ZNSs6resizeEyc _ZNSs6resizeEyc .text$_ZNSs6resizeEy _ZNSs6resizeEy .text$_ZNSs9push_backEc _ZNSs9push_backEc .text$_ZNSspLEc _ZNSspLEc .text$_ZNSs4_Rep7_M_grabERKSaIcES2_ _ZNSs4_Rep7_M_grabERKSaIcES2_ .text$_ZNSsC1ERKSs _ZNSsC1ERKSs .text$_ZNSsC2ERKSs _ZNSsC2ERKSs .text$_ZNSs6assignERKSs _ZNSs6assignERKSs .text$_ZNSsaSERKSs _ZNSsaSERKSs .text$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ .text$_ZStplIcSt11char_traits�      IcESaIcEESbIT_T0_T1_ES3_RKS6_ _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ES3_RKS6_ .text$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ .text$_ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag _ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag .text$_ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE _ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE .text$_ZNSsC1IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE _ZNSsC1IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE .text$_ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag _ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag .text$_ZNSsC2ERKSsyRKSaIcE _ZNSsC2ERKSsyRKSaIcE .text$_ZNSsC1ERKSsyRKSaIcE _ZNSsC1ERKSsyRKSaIcE .text$_ZNSsC2ERKSsyy _ZNSsC2ERKSsyy .text$_ZNSsC1ERKSsyy _ZNSsC1ERKSsyy .text$_ZNKSs6substrEyy _ZNKSs6substrEyy .text$_ZNSsC2ERKSsyyRKS�      aIcE _ZNSsC2ERKSsyyRKSaIcE .text$_ZNSsC1ERKSsyyRKSaIcE _ZNSsC1ERKSsyyRKSaIcE .text$_ZNSsC2IPcEET_S1_RKSaIcE _ZNSsC2IPcEET_S1_RKSaIcE .text$_ZNSsC1IPcEET_S1_RKSaIcE _ZNSsC1IPcEET_S1_RKSaIcE .text$_ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag _ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag .text$_ZNSsC2EPKcyRKSaIcE _ZNSsC2EPKcyRKSaIcE .text$_ZNSsC1EPKcyRKSaIcE _ZNSsC1EPKcyRKSaIcE .text$_ZNSs7replaceEyyPKcy _ZNSs7replaceEyyPKcy .text$_ZNSs7replaceEyyRKSs _ZNSs7replaceEyyRKSs .text$_ZNSs7replaceEyyRKSsyy _ZNSs7replaceEyyRKSsyy .text$_ZNSs7replaceEyyPKc _ZNSs7replaceEyyPKc .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcy _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcy .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc .text$_ZNSs7replaceEN9__gnu_cxx17__no�      rmal_iteratorIPcSsEES2_S1_S1_ _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S1_S1_ .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_St16initializer_listIcE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_St16initializer_listIcE .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ .text$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ .text$_ZNSsC2EPKcRKSaIcE _ZNSsC2EPKcRKSaIcE .text$_ZNSsC1EPKcRKSaIcE _ZNSsC1EPKcRKSaIcE .text$_ZNSsC2ESt16initializer_listIcERKSaIcE _ZNSsC2ESt16initializer_listIcERKSaIcE .text$_ZNSsC1ESt16initializer_listIcERKSaIcE _ZNSsC1ESt16initializer_listIcERKSaIcE .text$_ZNSsC2IPKcEET_S2_RKSaIcE _ZNSsC2IPKcEET_S2_RKSaIcE .text$_ZNSsC1IPKcEET_S2_RKSaIcE _ZNSsC1IPKcEET_�      S2_RKSaIcE .text$_ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ _ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ .text$_ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_T0_EES8_ _ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_T0_EES8_ _ZNSt13random_device7_M_initERKSs _ZNSt13random_device14_M_init_pretr1ERKSs .rdata$_ZNSs4_Rep11_S_terminalE .rdata$_ZNSs4_Rep11_S_max_sizeE .rdata$_ZNSs4nposE .xdata$_ZNKSs7_M_dataEv .pdata$_ZNKSs7_M_dataEv .xdata$_ZNSs7_M_dataEPc .pdata$_ZNSs7_M_dataEPc .xdata$_ZNKSs6_M_repEv .pdata$_ZNKSs6_M_repEv .xdata$_ZNKSs9_M_ibeginEv .pdata$_ZNKSs9_M_ibeginEv .xdata$_ZNKSs7_M_iendEv .pdata$_ZNKSs7_M_iendEv .xdata$_ZNKSs8_M_checkEyPKc .pdata$_ZNKSs8_M_checkEyPKc .xdata$_ZNKSs15_M_check_lengthEyyPKc .pdata$_ZNKSs15_M_check_lengthEyyPKc .xdata$_ZNKSs8_M_limitEyy .pdata$_ZNKSs8_M_limitEyy .xdata$_ZNKSs11_M_disjunctEPKc .pdata$_ZNKSs11_M_disjunctEPKc .xdata$_ZNSs7_M_copyEPcPKcy .pdata$_ZNSs7_M_copyEPcPKcy .xdata$_ZNSs7_M_moveEPcPKcy .pdata$_ZNSs7_M_moveEPcPKc�      y .xdata$_ZNSs9_M_assignEPcyc .pdata$_ZNSs9_M_assignEPcyc .xdata$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ .pdata$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ .xdata$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ .pdata$_ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ .xdata$_ZNSs13_S_copy_charsEPcS_S_ .pdata$_ZNSs13_S_copy_charsEPcS_S_ .xdata$_ZNSs13_S_copy_charsEPcPKcS1_ .pdata$_ZNSs13_S_copy_charsEPcPKcS1_ .xdata$_ZNSs10_S_compareEyy .pdata$_ZNSs10_S_compareEyy .xdata$_ZNSs12_S_empty_repEv .pdata$_ZNSs12_S_empty_repEv .xdata$_ZNSsD2Ev .pdata$_ZNSsD2Ev .xdata$_ZNSsD1Ev .pdata$_ZNSsD1Ev .xdata$_ZNKSs5beginEv .pdata$_ZNKSs5beginEv .xdata$_ZNKSs3endEv .pdata$_ZNKSs3endEv .xdata$_ZNKSs6rbeginEv .pdata$_ZNKSs6rbeginEv .xdata$_ZNKSs4rendEv .pdata$_ZNKSs4rendEv .xdata$_ZNKSs6cbeginEv .pdata$_ZNKSs6cbeginEv .xdata$_ZNKSs4cendEv .pdata$_ZNKSs4cendEv .xdata$_ZNKSs7crbeginEv .pdata$_ZNKSs7crbeginEv .xdata$_ZNKSs5crendEv .pdata$_ZNKSs5cr�      endEv .xdata$_ZNKSs4sizeEv .pdata$_ZNKSs4sizeEv .xdata$_ZNKSs6lengthEv .pdata$_ZNKSs6lengthEv .xdata$_ZNKSs8max_sizeEv .pdata$_ZNKSs8max_sizeEv .xdata$_ZNKSs8capacityEv .pdata$_ZNKSs8capacityEv .xdata$_ZNKSs5emptyEv .pdata$_ZNKSs5emptyEv .xdata$_ZNKSsixEy .pdata$_ZNKSsixEy .xdata$_ZNKSs2atEy .pdata$_ZNKSs2atEy .xdata$_ZNKSs5frontEv .pdata$_ZNKSs5frontEv .xdata$_ZNKSs4backEv .pdata$_ZNKSs4backEv .xdata$_ZNKSs4copyEPcyy .pdata$_ZNKSs4copyEPcyy .xdata$_ZNSs4swapERSs .pdata$_ZNSs4swapERSs .xdata$_ZNSsaSEOSs .pdata$_ZNSsaSEOSs .xdata$_ZNSs6assignEOSs .pdata$_ZNSs6assignEOSs .xdata$_ZNKSs5c_strEv .pdata$_ZNKSs5c_strEv .xdata$_ZNKSs4dataEv .pdata$_ZNKSs4dataEv .xdata$_ZNKSs13get_allocatorEv .pdata$_ZNKSs13get_allocatorEv .xdata$_ZNKSs4findEPKcyy .pdata$_ZNKSs4findEPKcyy .xdata$_ZNKSs4findERKSsy .pdata$_ZNKSs4findERKSsy .xdata$_ZNKSs4findEPKcy .pdata$_ZNKSs4findEPKcy .xdata$_ZNKSs4findEcy .pdata$_ZNKSs4findEcy .xdata$_ZNKSs5rfindEPKcyy .pdata$_ZNKSs5rfindEPKcyy .xdata$_ZNKSs5rfindERKSsy .pdata$_ZNKSs5rfindERK�      Ssy .xdata$_ZNKSs5rfindEPKcy .pdata$_ZNKSs5rfindEPKcy .xdata$_ZNKSs5rfindEcy .pdata$_ZNKSs5rfindEcy .xdata$_ZNKSs13find_first_ofEPKcyy .pdata$_ZNKSs13find_first_ofEPKcyy .xdata$_ZNKSs13find_first_ofERKSsy .pdata$_ZNKSs13find_first_ofERKSsy .xdata$_ZNKSs13find_first_ofEPKcy .pdata$_ZNKSs13find_first_ofEPKcy .xdata$_ZNKSs13find_first_ofEcy .pdata$_ZNKSs13find_first_ofEcy .xdata$_ZNKSs12find_last_ofEPKcyy .pdata$_ZNKSs12find_last_ofEPKcyy .xdata$_ZNKSs12find_last_ofERKSsy .pdata$_ZNKSs12find_last_ofERKSsy .xdata$_ZNKSs12find_last_ofEPKcy .pdata$_ZNKSs12find_last_ofEPKcy .xdata$_ZNKSs12find_last_ofEcy .pdata$_ZNKSs12find_last_ofEcy .xdata$_ZNKSs17find_first_not_ofEPKcyy .pdata$_ZNKSs17find_first_not_ofEPKcyy .xdata$_ZNKSs17find_first_not_ofERKSsy .pdata$_ZNKSs17find_first_not_ofERKSsy .xdata$_ZNKSs17find_first_not_ofEPKcy .pdata$_ZNKSs17find_first_not_ofEPKcy .xdata$_ZNKSs17find_first_not_ofEcy .pdata$_ZNKSs17find_first_not_ofEcy .xdata$_ZNKSs16find_last_not_ofEPKcyy .pdata$_ZNKSs16find_last_not_ofEPKcyy �      .xdata$_ZNKSs16find_last_not_ofERKSsy .pdata$_ZNKSs16find_last_not_ofERKSsy .xdata$_ZNKSs16find_last_not_ofEPKcy .pdata$_ZNKSs16find_last_not_ofEPKcy .xdata$_ZNKSs16find_last_not_ofEcy .pdata$_ZNKSs16find_last_not_ofEcy .xdata$_ZNKSs7compareERKSs .pdata$_ZNKSs7compareERKSs .xdata$_ZNKSs7compareEyyRKSs .pdata$_ZNKSs7compareEyyRKSs .xdata$_ZNKSs7compareEyyRKSsyy .pdata$_ZNKSs7compareEyyRKSsyy .xdata$_ZNKSs7compareEPKc .pdata$_ZNKSs7compareEPKc .xdata$_ZNKSs7compareEyyPKc .pdata$_ZNKSs7compareEyyPKc .xdata$_ZNKSs7compareEyyPKcy .pdata$_ZNKSs7compareEyyPKcy .xdata$_ZNSs12_Alloc_hiderC2EPcRKSaIcE .pdata$_ZNSs12_Alloc_hiderC2EPcRKSaIcE .xdata$_ZNSs12_Alloc_hiderC1EPcRKSaIcE .pdata$_ZNSs12_Alloc_hiderC1EPcRKSaIcE .xdata$_ZNSs4_Rep12_S_empty_repEv .pdata$_ZNSs4_Rep12_S_empty_repEv .xdata$_ZNKSs4_Rep12_M_is_leakedEv .pdata$_ZNKSs4_Rep12_M_is_leakedEv .xdata$_ZNKSs4_Rep12_M_is_sharedEv .pdata$_ZNKSs4_Rep12_M_is_sharedEv .xdata$_ZNSs4_Rep13_M_set_leakedEv .pdata$_ZNSs4_Rep13_M_set_leakedEv .xdata$_ZNSs4_Rep15_M_�      set_sharableEv .pdata$_ZNSs4_Rep15_M_set_sharableEv .xdata$_ZNSs4_Rep26_M_set_length_and_sharableEy .pdata$_ZNSs4_Rep26_M_set_length_and_sharableEy .xdata$_ZNSs4_Rep10_M_refdataEv .pdata$_ZNSs4_Rep10_M_refdataEv .xdata$_ZNSs4_Rep9_S_createEyyRKSaIcE .pdata$_ZNSs4_Rep9_S_createEyyRKSaIcE .xdata$_ZNSs9_M_mutateEyyy .pdata$_ZNSs9_M_mutateEyyy .xdata$_ZNSs12_M_leak_hardEv .pdata$_ZNSs12_M_leak_hardEv .xdata$_ZNSs7_M_leakEv .pdata$_ZNSs7_M_leakEv .xdata$_ZNSs4rendEv .pdata$_ZNSs4rendEv .xdata$_ZNSs5frontEv .pdata$_ZNSs5frontEv .xdata$_ZNSsixEy .pdata$_ZNSsixEy .xdata$_ZNSs5beginEv .pdata$_ZNSs5beginEv .xdata$_ZNSs6rbeginEv .pdata$_ZNSs6rbeginEv .xdata$_ZNSs3endEv .pdata$_ZNSs3endEv .xdata$_ZNSs4backEv .pdata$_ZNSs4backEv .xdata$_ZNSs2atEy .pdata$_ZNSs2atEy .xdata$_ZNSs5clearEv .pdata$_ZNSs5clearEv .xdata$_ZNSs5eraseEyy .pdata$_ZNSs5eraseEyy .xdata$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE .pdata$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE .xdata$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSs�      EES2_ .pdata$_ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEES2_ .xdata$_ZNSs14_M_replace_auxEyyyc .pdata$_ZNSs14_M_replace_auxEyyyc .xdata$_ZNSs6assignEyc .pdata$_ZNSs6assignEyc .xdata$_ZNSsaSEc .pdata$_ZNSsaSEc .xdata$_ZNSs6insertEyyc .pdata$_ZNSs6insertEyyc .xdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc .pdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc .xdata$_ZNSs7replaceEyyyc .pdata$_ZNSs7replaceEyyyc .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_yc .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_yc .xdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEyc .pdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEyc .xdata$_ZNSs15_M_replace_safeEyyPKcy .pdata$_ZNSs15_M_replace_safeEyyPKcy .xdata$_ZNSs6assignEPKcy .pdata$_ZNSs6assignEPKcy .xdata$_ZNSsaSESt16initializer_listIcE .pdata$_ZNSsaSESt16initializer_listIcE .xdata$_ZNSs6assignERKSsyy .pdata$_ZNSs6assignERKSsyy .xdata$_ZNSs6assignEPKc .pdata$_ZNSs6assignEPKc .xdata$_ZNSsaSEPKc .pdata$_ZNSsa�      SEPKc .xdata$_ZNSs6assignESt16initializer_listIcE .pdata$_ZNSs6assignESt16initializer_listIcE .xdata$_ZNSs6insertEyPKcy .pdata$_ZNSs6insertEyPKcy .xdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE .pdata$_ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE .xdata$_ZNSs6insertEyRKSsyy .pdata$_ZNSs6insertEyRKSsyy .xdata$_ZNSs6insertEyPKc .pdata$_ZNSs6insertEyPKc .xdata$_ZNSs6insertEyRKSs .pdata$_ZNSs6insertEyRKSs .xdata$_ZNSs8pop_backEv .pdata$_ZNSs8pop_backEv .xdata$_ZNSs12_S_constructEycRKSaIcE .pdata$_ZNSs12_S_constructEycRKSaIcE .xdata$_ZNSsC2Ev .pdata$_ZNSsC2Ev .xdata$_ZNSsC1Ev .pdata$_ZNSsC1Ev .xdata$_ZNSsC2ERKSaIcE .pdata$_ZNSsC2ERKSaIcE .xdata$_ZNSsC1ERKSaIcE .pdata$_ZNSsC1ERKSaIcE .xdata$_ZNSsC2EycRKSaIcE .pdata$_ZNSsC2EycRKSaIcE .xdata$_ZNSsC1EycRKSaIcE .pdata$_ZNSsC1EycRKSaIcE .xdata$_ZNSsC2EOSs .pdata$_ZNSsC2EOSs .xdata$_ZNSsC1EOSs .pdata$_ZNSsC1EOSs .xdata$_ZNSs18_S_construct_aux_2EycRKSaIcE .pdata$_ZNSs18_S_construct_aux_2EycRKSaIcE .xdata�      $_ZNSs4_Rep10_M_disposeERKSaIcE .pdata$_ZNSs4_Rep10_M_disposeERKSaIcE .xdata$_ZNSs4_Rep10_M_destroyERKSaIcE .pdata$_ZNSs4_Rep10_M_destroyERKSaIcE .xdata$_ZNSs4_Rep10_M_refcopyEv .pdata$_ZNSs4_Rep10_M_refcopyEv .xdata$_ZNSs4_Rep8_M_cloneERKSaIcEy .pdata$_ZNSs4_Rep8_M_cloneERKSaIcEy .xdata$_ZNSs7reserveEy .pdata$_ZNSs7reserveEy .xdata$_ZNSs13shrink_to_fitEv .pdata$_ZNSs13shrink_to_fitEv .xdata$_ZNSs6appendERKSs .pdata$_ZNSs6appendERKSs .xdata$_ZNSspLERKSs .pdata$_ZNSspLERKSs .xdata$_ZNSs6appendERKSsyy .pdata$_ZNSs6appendERKSsyy .xdata$_ZNSs6appendEPKcy .pdata$_ZNSs6appendEPKcy .xdata$_ZNSspLESt16initializer_listIcE .pdata$_ZNSspLESt16initializer_listIcE .xdata$_ZNSs6appendEPKc .pdata$_ZNSs6appendEPKc .xdata$_ZNSspLEPKc .pdata$_ZNSspLEPKc .xdata$_ZNSs6appendESt16initializer_listIcE .pdata$_ZNSs6appendESt16initializer_listIcE .text$_ZNSs6appendEyc.part.20 .xdata$_ZNSs6appendEyc.part.20 .pdata$_ZNSs6appendEyc.part.20 .xdata$_ZNSs6appendEyc .pdata$_ZNSs6appendEyc .xdata$_ZNSs6resizeEyc .pdata$_ZNSs6resizeEy�      c .xdata$_ZNSs6resizeEy .pdata$_ZNSs6resizeEy .xdata$_ZNSs9push_backEc .pdata$_ZNSs9push_backEc .xdata$_ZNSspLEc .pdata$_ZNSspLEc .xdata$_ZNSs4_Rep7_M_grabERKSaIcES2_ .pdata$_ZNSs4_Rep7_M_grabERKSaIcES2_ .xdata$_ZNSsC1ERKSs .pdata$_ZNSsC1ERKSs .xdata$_ZNSsC2ERKSs .pdata$_ZNSsC2ERKSs .xdata$_ZNSs6assignERKSs .pdata$_ZNSs6assignERKSs .xdata$_ZNSsaSERKSs .pdata$_ZNSsaSERKSs .xdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ .pdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ .xdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ES3_RKS6_ .pdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ES3_RKS6_ .xdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ .pdata$_ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ .xdata$_ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag .pdata$_ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag .xdata$_ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE�       .pdata$_ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE .xdata$_ZNSsC1IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE .pdata$_ZNSsC1IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE .xdata$_ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag .pdata$_ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag .xdata$_ZNSsC2ERKSsyRKSaIcE .pdata$_ZNSsC2ERKSsyRKSaIcE .xdata$_ZNSsC1ERKSsyRKSaIcE .pdata$_ZNSsC1ERKSsyRKSaIcE .xdata$_ZNSsC2ERKSsyy .pdata$_ZNSsC2ERKSsyy .xdata$_ZNSsC1ERKSsyy .pdata$_ZNSsC1ERKSsyy .xdata$_ZNKSs6substrEyy .pdata$_ZNKSs6substrEyy .xdata$_ZNSsC2ERKSsyyRKSaIcE .pdata$_ZNSsC2ERKSsyyRKSaIcE .xdata$_ZNSsC1ERKSsyyRKSaIcE .pdata$_ZNSsC1ERKSsyyRKSaIcE .xdata$_ZNSsC2IPcEET_S1_RKSaIcE .pdata$_ZNSsC2IPcEET_S1_RKSaIcE .xdata$_ZNSsC1IPcEET_S1_RKSaIcE .pdata$_ZNSsC1IPcEET_S1_RKSaIcE .xdata$_ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag .pdata$_ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag .xdata$_ZNSsC2EPKcyRKSaIcE .pdata$_ZNS�      sC2EPKcyRKSaIcE .xdata$_ZNSsC1EPKcyRKSaIcE .pdata$_ZNSsC1EPKcyRKSaIcE .xdata$_ZNSs7replaceEyyPKcy .pdata$_ZNSs7replaceEyyPKcy .xdata$_ZNSs7replaceEyyRKSs .pdata$_ZNSs7replaceEyyRKSs .xdata$_ZNSs7replaceEyyRKSsyy .pdata$_ZNSs7replaceEyyRKSsyy .xdata$_ZNSs7replaceEyyPKc .pdata$_ZNSs7replaceEyyPKc .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcy .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcy .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S1_S1_ .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S1_S1_ .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPc�      SsEES2_St16initializer_listIcE .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_St16initializer_listIcE .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ .xdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ .pdata$_ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ .xdata$_ZNSsC2EPKcRKSaIcE .pdata$_ZNSsC2EPKcRKSaIcE .xdata$_ZNSsC1EPKcRKSaIcE .pdata$_ZNSsC1EPKcRKSaIcE .xdata$_ZNSsC2ESt16initializer_listIcERKSaIcE .pdata$_ZNSsC2ESt16initializer_listIcERKSaIcE .xdata$_ZNSsC1ESt16initializer_listIcERKSaIcE .pdata$_ZNSsC1ESt16initializer_listIcERKSaIcE .xdata$_ZNSsC2IPKcEET_S2_RKSaIcE .pdata$_ZNSsC2IPKcEET_S2_RKSaIcE .xdata$_ZNSsC1IPKcEET_S2_RKSaIcE .pdata$_ZNSsC1IPKcEET_S2_RKSaIcE .xdata$_ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ .pdata$_ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ .xdata$_ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_�      T0_EES8_ .pdata$_ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_T0_EES8_ .text$_ZNSt13random_device7_M_initERKSs .xdata$_ZNSt13random_device7_M_initERKSs .pdata$_ZNSt13random_device7_M_initERKSs .text$_ZNSt13random_device14_M_init_pretr1ERKSs .xdata$_ZNSt13random_device14_M_init_pretr1ERKSs .pdata$_ZNSt13random_device14_M_init_pretr1ERKSs .text$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_dataEv _ZNKSbIwSt11char_traitsIwESaIwEE7_M_dataEv .text$_ZNSbIwSt11char_traitsIwESaIwEE7_M_dataEPw _ZNSbIwSt11char_traitsIwESaIwEE7_M_dataEPw .text$_ZNKSbIwSt11char_traitsIwESaIwEE6_M_repEv _ZNKSbIwSt11char_traitsIwESaIwEE6_M_repEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE9_M_ibeginEv _ZNKSbIwSt11char_traitsIwESaIwEE9_M_ibeginEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_iendEv _ZNKSbIwSt11char_traitsIwESaIwEE7_M_iendEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_checkEyPKc _ZNKSbIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .text$_ZNKSbIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc _ZNKSbIwSt11char_traitsIwESaIwEE15_M_check_lengt�      hEyyPKc .text$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_limitEyy _ZNKSbIwSt11char_traitsIwESaIwEE8_M_limitEyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw _ZNKSbIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .text$_ZNSbIwSt11char_traitsIwESaIwEE7_M_copyEPwPKwy _ZNSbIwSt11char_traitsIwESaIwEE7_M_copyEPwPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE7_M_moveEPwPKwy _ZNSbIwSt11char_traitsIwESaIwEE7_M_moveEPwPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE9_M_assignEPwyw _ZNSbIwSt11char_traitsIwESaIwEE9_M_assignEPwyw .text$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS3_S2_EES6_ _ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS3_S2_EES6_ .text$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS2_EES8_ _ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS2_EES8_ .text$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS3_S3_ _ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS3_S3_ .text$_Z�      NSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS5_ _ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS5_ .text$_ZNSbIwSt11char_traitsIwESaIwEE10_S_compareEyy _ZNSbIwSt11char_traitsIwESaIwEE10_S_compareEyy .text$_ZNSbIwSt11char_traitsIwESaIwEE12_S_empty_repEv _ZNSbIwSt11char_traitsIwESaIwEE12_S_empty_repEv .data$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep20_S_empty_rep_storageE .text$_ZNSbIwSt11char_traitsIwESaIwEED2Ev _ZNSbIwSt11char_traitsIwESaIwEED2Ev .text$_ZNSbIwSt11char_traitsIwESaIwEED1Ev _ZNSbIwSt11char_traitsIwESaIwEED1Ev .text$_ZNKSbIwSt11char_traitsIwESaIwEE5beginEv _ZNKSbIwSt11char_traitsIwESaIwEE5beginEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE3endEv _ZNKSbIwSt11char_traitsIwESaIwEE3endEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE6rbeginEv _ZNKSbIwSt11char_traitsIwESaIwEE6rbeginEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4rendEv _ZNKSbIwSt11char_traitsIwESaIwEE4rendEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE6cbeginEv _ZNKSbIwSt11char_traitsIwESaIwEE6cbeginEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4cendE�      v _ZNKSbIwSt11char_traitsIwESaIwEE4cendEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE7crbeginEv _ZNKSbIwSt11char_traitsIwESaIwEE7crbeginEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE5crendEv _ZNKSbIwSt11char_traitsIwESaIwEE5crendEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4sizeEv _ZNKSbIwSt11char_traitsIwESaIwEE4sizeEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE6lengthEv _ZNKSbIwSt11char_traitsIwESaIwEE6lengthEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE8max_sizeEv _ZNKSbIwSt11char_traitsIwESaIwEE8max_sizeEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE8capacityEv _ZNKSbIwSt11char_traitsIwESaIwEE8capacityEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE5emptyEv _ZNKSbIwSt11char_traitsIwESaIwEE5emptyEv .text$_ZNKSbIwSt11char_traitsIwESaIwEEixEy _ZNKSbIwSt11char_traitsIwESaIwEEixEy .text$_ZNKSbIwSt11char_traitsIwESaIwEE2atEy _ZNKSbIwSt11char_traitsIwESaIwEE2atEy .text$_ZNKSbIwSt11char_traitsIwESaIwEE5frontEv _ZNKSbIwSt11char_traitsIwESaIwEE5frontEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4backEv _ZNKSbIwSt11char_traitsIwESaIwEE4backEv .text$�      _ZNKSbIwSt11char_traitsIwESaIwEE4copyEPwyy _ZNKSbIwSt11char_traitsIwESaIwEE4copyEPwyy .text$_ZNSbIwSt11char_traitsIwESaIwEE4swapERS2_ _ZNSbIwSt11char_traitsIwESaIwEE4swapERS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEEaSEOS2_ _ZNSbIwSt11char_traitsIwESaIwEEaSEOS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignEOS2_ _ZNSbIwSt11char_traitsIwESaIwEE6assignEOS2_ .text$_ZNKSbIwSt11char_traitsIwESaIwEE5c_strEv _ZNKSbIwSt11char_traitsIwESaIwEE5c_strEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4dataEv _ZNKSbIwSt11char_traitsIwESaIwEE4dataEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE13get_allocatorEv _ZNKSbIwSt11char_traitsIwESaIwEE13get_allocatorEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE4findERKS2_y _ZNKSbIwSt11char_traitsIwESaIwEE4findERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE4findEwy _ZNKSbIwSt11char_traitsIwESaIwEE4findEwy .text$_ZNKSb�      IwSt11char_traitsIwESaIwEE5rfindEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindERKS2_y _ZNKSbIwSt11char_traitsIwESaIwEE5rfindERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEwy _ZNKSbIwSt11char_traitsIwESaIwEE5rfindEwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofERKS2_y _ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEwy _ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofERKS2_y _ZNKSbIwSt11char_traitsIwESa�      IwEE12find_last_ofERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEwy _ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS2_y _ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy _ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy _ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .text$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS2_y _ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS2_y .text$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_�      not_ofEPKwy _ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy _ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareERKS2_ _ZNKSbIwSt11char_traitsIwESaIwEE7compareERKS2_ .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_ _ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_ .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_yy _ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_yy .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEPKw _ZNKSbIwSt11char_traitsIwESaIwEE7compareEPKw .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKw _ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKw .text$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKwy _ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS1_ _ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS1_ _ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hide�      rC1EPwRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep12_S_empty_repEv _ZNSbIwSt11char_traitsIwESaIwEE4_Rep12_S_empty_repEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_leakedEv _ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_leakedEv .text$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_sharedEv _ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_sharedEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep13_M_set_leakedEv _ZNSbIwSt11char_traitsIwESaIwEE4_Rep13_M_set_leakedEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep15_M_set_sharableEv _ZNSbIwSt11char_traitsIwESaIwEE4_Rep15_M_set_sharableEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep26_M_set_length_and_sharableEy _ZNSbIwSt11char_traitsIwESaIwEE4_Rep26_M_set_length_and_sharableEy .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refdataEv _ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refdataEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep9_S_createEyyRKS1_ _ZNSbIwSt11char_traitsIwESaIwEE4_Rep9_S_createEyyRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE9_M_mutateEyyy _ZNSbIwSt11char_�      traitsIwESaIwEE9_M_mutateEyyy .text$_ZNSbIwSt11char_traitsIwESaIwEE12_M_leak_hardEv _ZNSbIwSt11char_traitsIwESaIwEE12_M_leak_hardEv .text$_ZNSbIwSt11char_traitsIwESaIwEE7_M_leakEv _ZNSbIwSt11char_traitsIwESaIwEE7_M_leakEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4rendEv _ZNSbIwSt11char_traitsIwESaIwEE4rendEv .text$_ZNSbIwSt11char_traitsIwESaIwEE5frontEv _ZNSbIwSt11char_traitsIwESaIwEE5frontEv .text$_ZNSbIwSt11char_traitsIwESaIwEE5beginEv _ZNSbIwSt11char_traitsIwESaIwEE5beginEv .text$_ZNSbIwSt11char_traitsIwESaIwEEixEy _ZNSbIwSt11char_traitsIwESaIwEEixEy .text$_ZNSbIwSt11char_traitsIwESaIwEE6rbeginEv _ZNSbIwSt11char_traitsIwESaIwEE6rbeginEv .text$_ZNSbIwSt11char_traitsIwESaIwEE4backEv _ZNSbIwSt11char_traitsIwESaIwEE4backEv .text$_ZNSbIwSt11char_traitsIwESaIwEE3endEv _ZNSbIwSt11char_traitsIwESaIwEE3endEv .text$_ZNSbIwSt11char_traitsIwESaIwEE2atEy _ZNSbIwSt11char_traitsIwESaIwEE2atEy .text$_ZNSbIwSt11char_traitsIwESaIwEE5clearEv _ZNSbIwSt11char_traitsIwESaIwEE5clearEv .text$_ZNSbIwSt11char_traitsIwESaIwEE5er�      aseEyy _ZNSbIwSt11char_traitsIwESaIwEE5eraseEyy .text$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EE _ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EE .text$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_ _ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_ .text$_ZNSbIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw _ZNSbIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignEyw _ZNSbIwSt11char_traitsIwESaIwEE6assignEyw .text$_ZNSbIwSt11char_traitsIwESaIwEEaSEw _ZNSbIwSt11char_traitsIwESaIwEEaSEw .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyyw _ZNSbIwSt11char_traitsIwESaIwEE6insertEyyw .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEw _ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEw .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyyw _ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyyw .text$_ZNS�      bIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_yw _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_yw .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEyw _ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEyw .text$_ZNSbIwSt11char_traitsIwESaIwEE15_M_replace_safeEyyPKwy _ZNSbIwSt11char_traitsIwESaIwEE15_M_replace_safeEyyPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKwy _ZNSbIwSt11char_traitsIwESaIwEE6assignEPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE _ZNSbIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_yy _ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_yy .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKw _ZNSbIwSt11char_traitsIwESaIwEE6assignEPKw .text$_ZNSbIwSt11char_traitsIwESaIwEEaSEPKw _ZNSbIwSt11char_traitsIwESaIwEEaSEPKw .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE _ZNSbIwSt�      11char_traitsIwESaIwEE6assignESt16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKwy _ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EESt16initializer_listIwE _ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EESt16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_yy _ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_yy .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKw _ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKw .text$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_ _ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE8pop_backEv _ZNSbIwSt11char_traitsIwESaIwEE8pop_backEv .text$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructEywRKS1_ _ZNSbIwSt11char_traitsIwESaIwEE12_S_constructEywRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2EywRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2EywRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1EywRKS1_ _ZNSbIwSt11char_trai�      tsIwESaIwEEC1EywRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE18_S_construct_aux_2EywRKS1_ _ZNSbIwSt11char_traitsIwESaIwEE18_S_construct_aux_2EywRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2Ev _ZNSbIwSt11char_traitsIwESaIwEEC2Ev .text$_ZNSbIwSt11char_traitsIwESaIwEEC1Ev _ZNSbIwSt11char_traitsIwESaIwEEC1Ev .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2ERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1ERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2EOS2_ _ZNSbIwSt11char_traitsIwESaIwEEC2EOS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1EOS2_ _ZNSbIwSt11char_traitsIwESaIwEEC1EOS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_disposeERKS1_ _ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_disposeERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_destroyERKS1_ _ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_destroyERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refcopyEv _ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refcopyEv .text$_ZNSbIwSt11char_traitsIwES�      aIwEE4_Rep8_M_cloneERKS1_y _ZNSbIwSt11char_traitsIwESaIwEE4_Rep8_M_cloneERKS1_y .text$_ZNSbIwSt11char_traitsIwESaIwEE7reserveEy _ZNSbIwSt11char_traitsIwESaIwEE7reserveEy .text$_ZNSbIwSt11char_traitsIwESaIwEE13shrink_to_fitEv _ZNSbIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_ _ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEEpLERKS2_ _ZNSbIwSt11char_traitsIwESaIwEEpLERKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_yy _ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_yy .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKwy _ZNSbIwSt11char_traitsIwESaIwEE6appendEPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE _ZNSbIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKw _ZNSbIwSt11char_traitsIwESaIwEE6appendEPKw .text$_ZNSbIwSt11char_traitsIwESaIwEEpLEPKw _ZNSbIwSt11char_traitsIwESaIwEEpLEPKw .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE _�      ZNSbIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE _ZNSbIwSt11char_traitsIwESaIwEE6appendEyw.part.25 .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw _ZNSbIwSt11char_traitsIwESaIwEE6appendEyw .text$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEyw _ZNSbIwSt11char_traitsIwESaIwEE6resizeEyw .text$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEy _ZNSbIwSt11char_traitsIwESaIwEE6resizeEy .text$_ZNSbIwSt11char_traitsIwESaIwEE9push_backEw _ZNSbIwSt11char_traitsIwESaIwEE9push_backEw .text$_ZNSbIwSt11char_traitsIwESaIwEEpLEw _ZNSbIwSt11char_traitsIwESaIwEEpLEw .text$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep7_M_grabERKS1_S5_ _ZNSbIwSt11char_traitsIwESaIwEE4_Rep7_M_grabERKS1_S5_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_ _ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_ _ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_ _ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEEaSERKS2_ _ZNSbIwSt11char_traitsIwESaIwEEaSERK�      S2_ .text$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_EPKS3_RKS6_ _ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_EPKS3_RKS6_ .text$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ES3_RKS6_ _ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ES3_RKS6_ .text$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ERKS6_S8_ _ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ERKS6_S8_ .text$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIN9__gnu_cxx17__normal_iteratorIPwS2_EEEES6_T_S8_RKS1_St20forward_iterator_tag _ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIN9__gnu_cxx17__normal_iteratorIPwS2_EEEES6_T_S8_RKS1_St20forward_iterator_tag .text$_ZNSbIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPwEES4_T_S5_RK�      S1_St20forward_iterator_tag _ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPwEES4_T_S5_RKS1_St20forward_iterator_tag .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yy _ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yy .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yy _ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yy .text$_ZNKSbIwSt11char_traitsIwESaIwEE6substrEyy _ZNKSbIwSt11char_traitsIwESaIwEE6substrEyy .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yyRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yyRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yyRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yyRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2IPwEET_S5_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2IPwEET_S5_RKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1IPwEET_S5_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1IPwEET_S5_RKS1_ .text$_ZNSbIwSt11char_tr�      aitsIwESaIwEE12_S_constructIPKwEEPwT_S7_RKS1_St20forward_iterator_tag _ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPKwEEPwT_S7_RKS1_St20forward_iterator_tag .text$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwyRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2EPKwyRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwyRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1EPKwyRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKwy _ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_yy _ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_yy .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKw _ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKw .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwy _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwy .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6�      _RKS2_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_RKS2_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKw _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKw .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S5_S5_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S5_S5_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwS8_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwS8_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_St16initializer_listIwE _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_St16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S6_S6_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIP�      wS2_EES6_S6_S6_ .text$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_NS4_IPKwS2_EES9_ _ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_NS4_IPKwS2_EES9_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2EPKwRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwRKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1EPKwRKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC2IPKwEET_S6_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC2IPKwEET_S6_RKS1_ .text$_ZNSbIwSt11char_traitsIwESaIwEEC1IPKwEET_S6_RKS1_ _ZNSbIwSt11char_traitsIwESaIwEEC1IPKwEET_S6_RKS1_ .text$_ZN9__gnu_cxxeqIPwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESB_ _ZN9__gnu_cxxeqIPwSbIwSt11char_traitsIwESaIwEEE�      EbRKNS_17__normal_iteratorIT_T0_EESB_ .text$_ZN9__gnu_cxxeqIPKwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESC_ _ZN9__gnu_cxxeqIPKwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESC_ .rdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep11_S_terminalE .rdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep11_S_max_sizeE .rdata$_ZNSbIwSt11char_traitsIwESaIwEE4nposE .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_dataEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_dataEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_dataEPw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_dataEPw .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE6_M_repEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE6_M_repEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE9_M_ibeginEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE9_M_ibeginEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_iendEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7_M_iendEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .xdata$_ZNKSbIwSt11char_trait�      sIwESaIwEE15_M_check_lengthEyyPKc .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_limitEyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE8_M_limitEyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_copyEPwPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_copyEPwPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_moveEPwPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_moveEPwPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE9_M_assignEPwyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE9_M_assignEPwyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS3_S2_EES6_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS3_S2_EES6_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS2_EES8_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_it�      eratorIPKwS2_EES8_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS3_S3_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS3_S3_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS5_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS5_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE10_S_compareEyy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE10_S_compareEyy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_empty_repEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_empty_repEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEED2Ev .pdata$_ZNSbIwSt11char_traitsIwESaIwEED2Ev .xdata$_ZNSbIwSt11char_traitsIwESaIwEED1Ev .pdata$_ZNSbIwSt11char_traitsIwESaIwEED1Ev .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5beginEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5beginEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE3endEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE3endEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE6rbeginEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE6rbeginEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4rendEv .pdata$_ZNKSbIwSt11cha�      r_traitsIwESaIwEE4rendEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE6cbeginEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE6cbeginEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4cendEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4cendEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7crbeginEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7crbeginEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5crendEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5crendEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4sizeEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4sizeEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE6lengthEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE6lengthEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE8max_sizeEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE8max_sizeEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE8capacityEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE8capacityEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5emptyEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5emptyEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEEixEy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEEixEy .xdata$_ZNKSbIwSt11char�      _traitsIwESaIwEE2atEy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE2atEy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5frontEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5frontEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4backEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4backEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4copyEPwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4copyEPwyy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4swapERS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4swapERS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEOS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEOS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEOS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEOS2_ .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5c_strEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5c_strEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4dataEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4dataEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE13get_allocatorEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE13get_allocatorEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwyy .pdata$_ZNKS�      bIwSt11char_traitsIwESaIwEE4findEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findERKS2_y .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4findEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindERKS2_y .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE5rfindEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofERKS2_y .xdata$_ZNKSbIwSt11ch�      ar_traitsIwESaIwEE13find_first_ofEPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE13find_first_ofEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofERKS2_y .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE12find_last_ofEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS2_y .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .�      pdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS2_y .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS2_y .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareERKS2_ .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareERKS2_ .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_ .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_ .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyRKS2_yy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compa�      reEyyRKS2_yy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEPKw .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEPKw .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKw .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKw .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKwy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE7compareEyyPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep12_S_empty_repEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep12_S_empty_repEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_leakedEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_leakedEv .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_sharedEv .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE4_Rep12_M_is_sharedEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep13_M_set_leakedEv .pda�      ta$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep13_M_set_leakedEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep15_M_set_sharableEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep15_M_set_sharableEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep26_M_set_length_and_sharableEy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep26_M_set_length_and_sharableEy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refdataEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refdataEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep9_S_createEyyRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep9_S_createEyyRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE9_M_mutateEyyy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE9_M_mutateEyyy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_M_leak_hardEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_M_leak_hardEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_leakEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7_M_leakEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4rendEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4rendEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5�      frontEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5frontEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5beginEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5beginEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEEixEy .pdata$_ZNSbIwSt11char_traitsIwESaIwEEixEy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6rbeginEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6rbeginEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4backEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4backEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE3endEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE3endEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE2atEy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE2atEy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5clearEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5clearEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEyy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEyy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EE .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx1�      7__normal_iteratorIPwS2_EES6_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEw .pdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_yw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_yw .xdata$_ZNSbIwSt11char_traitsIwESaIwE�      E6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EEyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE15_M_replace_safeEyyPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE15_M_replace_safeEyyPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_yy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignEPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEPKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEEaSEPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKwy .pdata$_ZNSbIwSt11char_traitsIw�      ESaIwEE6insertEyPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EESt16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS2_EESt16initializer_listIwE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_yy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6insertEyRKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE8pop_backEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE8pop_backEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructEywRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructEywRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EywRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EywRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EywRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EywRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE18_S_�      construct_aux_2EywRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE18_S_construct_aux_2EywRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2Ev .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2Ev .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1Ev .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1Ev .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EOS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EOS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EOS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EOS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_disposeERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_disposeERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_destroyERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_destroyERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refcopyEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep10_M_refcopyEv .xdata$_ZNSbIwSt1�      1char_traitsIwESaIwEE4_Rep8_M_cloneERKS1_y .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep8_M_cloneERKS1_y .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7reserveEy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7reserveEy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .pdata$_ZNSbIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEpLERKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEpLERKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendERKS2_yy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEEpLEPKw .pdata$_ZNSbIwSt11ch�      ar_traitsIwESaIwEEpLEPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE .text$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw.part.25 .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw.part.25 .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw.part.25 .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6appendEyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEyw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEyw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6resizeEy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE9push_backEw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE9push_backEw .xdata$_ZNSbIwSt11char_traitsIwESaIwEEpLEw .pdata$_ZNSbIwSt11char_traitsIwESaIwEEpLEw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep7_M_grabERKS1_S5_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE4_Rep7_M_grabERKS1_S5_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_ .pdata$_ZNSbIwSt11char_traitsIwE�      SaIwEEC1ERKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE6assignERKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEaSERKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEaSERKS2_ .xdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_EPKS3_RKS6_ .pdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_EPKS3_RKS6_ .xdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ES3_RKS6_ .pdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ES3_RKS6_ .xdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ERKS6_S8_ .pdata$_ZStplIwSt11char_traitsIwESaIwEESbIT_T0_T1_ERKS6_S8_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIN9__gnu_cxx17__normal_iteratorIPwS2_EEEES6_T_S8_RKS1_St20forward_iterator_tag .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIN9__gnu_cxx17__normal_iteratorIPwS2_EEEES6_T_S8_RKS1_St20forward_iterator_tag .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_�      S8_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS2_EEEET_S8_RKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPwEES4_T_S5_RKS1_St20forward_iterator_tag .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPwEES4_T_S5_RKS1_St20forward_iterator_tag .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yy .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yy .xdata$_ZNKSbIwSt11char_traitsIwESaIwEE6substrEyy .pdata$_ZNKSbIwSt11char_traitsIwESaIwEE6substrEyy .xdata$_ZNSbIwSt11char_traitsIwES�      aIwEEC2ERKS2_yyRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ERKS2_yyRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yyRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ERKS2_yyRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IPwEET_S5_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IPwEET_S5_RKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IPwEET_S5_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IPwEET_S5_RKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPKwEEPwT_S7_RKS1_St20forward_iterator_tag .pdata$_ZNSbIwSt11char_traitsIwESaIwEE12_S_constructIPKwEEPwT_S7_RKS1_St20forward_iterator_tag .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwyRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwyRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwyRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwyRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS�      2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_yy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyRKS2_yy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEyyPKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwy .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwy .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_RKS2_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_RKS2_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKw .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKw .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S5_S5_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S5_S5_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replac�      eEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwS8_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_PKwS8_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_St16initializer_listIwE .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_St16initializer_listIwE .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S6_S6_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_S6_S6_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_NS4_IPKwS2_EES9_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS2_EES6_NS4_IPKwS2_EES9_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2EPKwRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwRKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1EPKwRKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ESt16in�      itializer_listIwERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IPKwEET_S6_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC2IPKwEET_S6_RKS1_ .xdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IPKwEET_S6_RKS1_ .pdata$_ZNSbIwSt11char_traitsIwESaIwEEC1IPKwEET_S6_RKS1_ .xdata$_ZN9__gnu_cxxeqIPwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESB_ .pdata$_ZN9__gnu_cxxeqIPwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESB_ .xdata$_ZN9__gnu_cxxeqIPKwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESC_ .pdata$_ZN9__gnu_cxxeqIPKwSbIwSt11char_traitsIwESaIwEEEEbRKNS_17__normal_iteratorIT_T0_EESC_ .text$_ZNKSt5ctypeIcE8do_widenEc _ZNKSt5ctypeIcE8do_widenEc .text$_ZNKSt5ctypeIcE9do_narrowEcc _ZNKSt5ctypeIcE9do_narrowEcc _ZNSt5ctypeIcED2Ev .rdata$_ZTVSt5ctypeIcE _ZNSt5ctypeIcED1Ev �      _ZNSt5ctypeIwED2Ev .rdata$_ZTVSt5ctypeIwE .rdata$.refptr._ZTVSt21__ctype_abstract_baseIwE _ZNSt5ctypeIwED1Ev _ZNSt12ctype_bynameIwED2Ev _ZNSt12ctype_bynameIwED1Ev _ZNSt5ctypeIcED0Ev _ZNSt5ctypeIwED0Ev _ZNSt12ctype_bynameIwED0Ev .text$_ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc _ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc .text$_ZNKSt5ctypeIcE8do_widenEPKcS2_Pc _ZNKSt5ctypeIcE8do_widenEPKcS2_Pc _ZNKSt5ctypeIcE14_M_narrow_initEv _ZNKSt5ctypeIcE13_M_widen_initEv _ZNSt5ctypeIwEC2Ey _ZNSt5ctypeIwEC1Ey _ZNSt5ctypeIwEC2EPiy _ZNSt5ctypeIwEC1EPiy _ZNSt12ctype_bynameIwEC2EPKcy .rdata$_ZTVSt12ctype_bynameIwE _ZNSt12ctype_bynameIwEC1EPKcy .rdata$_ZTSSt10ctype_base .rdata$_ZTISt10ctype_base .rdata$_ZTSSt5ctypeIcE .rdata$_ZTISt5ctypeIcE .rdata$_ZTSSt21__ctype_abstract_baseIwE .rdata$_ZTISt21__ctype_abstract_baseIwE .rdata$_ZTSSt5ctypeIwE .rdata$_ZTISt5ctypeIwE .rdata$_ZTSSt12ctype_bynameIwE .rdata$_ZTISt12ctype_bynameIwE .xdata$_ZNKSt5ctypeIcE8do_widenEc .pdata$_ZNKSt5ctypeIcE8do_widenEc .xdata$_ZNKSt5ctypeIcE9do_narrowEcc .pdata$_�      ZNKSt5ctypeIcE9do_narrowEcc .text$_ZNSt5ctypeIcED2Ev .xdata$_ZNSt5ctypeIcED2Ev .pdata$_ZNSt5ctypeIcED2Ev .text$_ZNSt5ctypeIwED2Ev .xdata$_ZNSt5ctypeIwED2Ev .pdata$_ZNSt5ctypeIwED2Ev .text$_ZNSt12ctype_bynameIwED2Ev .xdata$_ZNSt12ctype_bynameIwED2Ev .pdata$_ZNSt12ctype_bynameIwED2Ev .text$_ZNSt5ctypeIcED0Ev .xdata$_ZNSt5ctypeIcED0Ev .pdata$_ZNSt5ctypeIcED0Ev .text$_ZNSt5ctypeIwED0Ev .xdata$_ZNSt5ctypeIwED0Ev .pdata$_ZNSt5ctypeIwED0Ev .text$_ZNSt12ctype_bynameIwED0Ev .xdata$_ZNSt12ctype_bynameIwED0Ev .pdata$_ZNSt12ctype_bynameIwED0Ev .xdata$_ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc .pdata$_ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc .xdata$_ZNKSt5ctypeIcE8do_widenEPKcS2_Pc .pdata$_ZNKSt5ctypeIcE8do_widenEPKcS2_Pc .text$_ZNKSt5ctypeIcE14_M_narrow_initEv .xdata$_ZNKSt5ctypeIcE14_M_narrow_initEv .pdata$_ZNKSt5ctypeIcE14_M_narrow_initEv .text$_ZNKSt5ctypeIcE13_M_widen_initEv .xdata$_ZNKSt5ctypeIcE13_M_widen_initEv .pdata$_ZNKSt5ctypeIcE13_M_widen_initEv .text$_ZNSt5ctypeIwEC2Ey .xdata$_ZNSt5ctypeIwEC2Ey .pdata$_ZNSt5ctype�      IwEC2Ey .text$_ZNSt5ctypeIwEC2EPiy .xdata$_ZNSt5ctypeIwEC2EPiy .pdata$_ZNSt5ctypeIwEC2EPiy .text$_ZNSt12ctype_bynameIwEC2EPKcy .xdata$_ZNSt12ctype_bynameIwEC2EPKcy .pdata$_ZNSt12ctype_bynameIwEC2EPKcy .rdata$_ZNSt5ctypeIcE10table_sizeE .data$_ZNSt5ctypeIwE2idE .data$_ZNSt5ctypeIcE2idE .rdata$_ZNSt10ctype_base5blankE .rdata$_ZNSt10ctype_base5graphE .rdata$_ZNSt10ctype_base5alnumE .rdata$_ZNSt10ctype_base6xdigitE .rdata$_ZNSt10ctype_base5punctE .rdata$_ZNSt10ctype_base5digitE .rdata$_ZNSt10ctype_base5alphaE .rdata$_ZNSt10ctype_base5lowerE .rdata$_ZNSt10ctype_base5upperE .rdata$_ZNSt10ctype_base5cntrlE .rdata$_ZNSt10ctype_base5printE .rdata$_ZNSt10ctype_base5spaceE _ZNKSt5ctypeIcE10do_toupperEc _ZNKSt5ctypeIcE10do_tolowerEc _ZNSt5ctypeIcE13classic_tableEv _ZZNSt5ctypeIcE13classic_tableEvE16_S_classic_table _ZNSt5ctypeIcEC2EPiPKtby .rdata$.refptr._ZTVSt5ctypeIcE _ZNSt5ctypeIcEC1EPiPKtby _ZNSt5ctypeIcEC2EPKtby _ZNSt5ctypeIcEC1EPKtby _ZNKSt5ctypeIcE10do_toupperEPcPKc _ZNKSt5ctypeIcE10do_tolowerEPcPKc .text$�      _ZNKSt5ctypeIcE10do_toupperEc .xdata$_ZNKSt5ctypeIcE10do_toupperEc .pdata$_ZNKSt5ctypeIcE10do_toupperEc .text$_ZNKSt5ctypeIcE10do_tolowerEc .xdata$_ZNKSt5ctypeIcE10do_tolowerEc .pdata$_ZNKSt5ctypeIcE10do_tolowerEc .text$_ZNSt5ctypeIcE13classic_tableEv .xdata$_ZNSt5ctypeIcE13classic_tableEv .pdata$_ZNSt5ctypeIcE13classic_tableEv .text$_ZNSt5ctypeIcEC2EPiPKtby .xdata$_ZNSt5ctypeIcEC2EPiPKtby .pdata$_ZNSt5ctypeIcEC2EPiPKtby .text$_ZNSt5ctypeIcEC2EPKtby .xdata$_ZNSt5ctypeIcEC2EPKtby .pdata$_ZNSt5ctypeIcEC2EPKtby .text$_ZNKSt5ctypeIcE10do_toupperEPcPKc .xdata$_ZNKSt5ctypeIcE10do_toupperEPcPKc .pdata$_ZNKSt5ctypeIcE10do_toupperEPcPKc .text$_ZNKSt5ctypeIcE10do_tolowerEPcPKc .xdata$_ZNKSt5ctypeIcE10do_tolowerEPcPKc .pdata$_ZNKSt5ctypeIcE10do_tolowerEPcPKc .rdata$_ZZNSt5ctypeIcE13classic_tableEvE16_S_classic_table _ZNSt12ctype_bynameIcED2Ev .rdata$_ZTVSt12ctype_bynameIcE _ZNSt12ctype_bynameIcED1Ev _ZNSt12ctype_bynameIcED0Ev _ZNSt12ctype_bynameIcEC2EPKcy _ZNSt12ctype_bynameIcEC1EPKcy _ZNKSt5ctypeIwE19_M_convert�      _to_wmaskEt _ZNKSt5ctypeIwE10do_toupperEw _ZNKSt5ctypeIwE10do_toupperEPwPKw _ZNKSt5ctypeIwE10do_tolowerEw _ZNKSt5ctypeIwE10do_tolowerEPwPKw _ZNKSt5ctypeIwE5do_isEtw _ZNKSt5ctypeIwE5do_isEPKwS2_Pt _ZNKSt5ctypeIwE10do_scan_isEtPKwS2_ _ZNKSt5ctypeIwE11do_scan_notEtPKwS2_ _ZNKSt5ctypeIwE8do_widenEc _ZNKSt5ctypeIwE8do_widenEPKcS2_Pw _ZNKSt5ctypeIwE9do_narrowEwc _ZNKSt5ctypeIwE9do_narrowEPKwS2_cPc _ZNSt5ctypeIwE19_M_initialize_ctypeEv .rdata$_ZTSSt12ctype_bynameIcE .rdata$_ZTISt12ctype_bynameIcE .text$_ZNSt12ctype_bynameIcED2Ev .xdata$_ZNSt12ctype_bynameIcED2Ev .pdata$_ZNSt12ctype_bynameIcED2Ev .text$_ZNSt12ctype_bynameIcED0Ev .xdata$_ZNSt12ctype_bynameIcED0Ev .pdata$_ZNSt12ctype_bynameIcED0Ev .text$_ZNSt12ctype_bynameIcEC2EPKcy .xdata$_ZNSt12ctype_bynameIcEC2EPKcy .pdata$_ZNSt12ctype_bynameIcEC2EPKcy .text$_ZNKSt5ctypeIwE19_M_convert_to_wmaskEt .xdata$_ZNKSt5ctypeIwE19_M_convert_to_wmaskEt .pdata$_ZNKSt5ctypeIwE19_M_convert_to_wmaskEt .text$_ZNKSt5ctypeIwE10do_toupperEw .xdata$_ZNKSt5ctypeIwE10do_toupperEw�       .pdata$_ZNKSt5ctypeIwE10do_toupperEw .text$_ZNKSt5ctypeIwE10do_toupperEPwPKw .xdata$_ZNKSt5ctypeIwE10do_toupperEPwPKw .pdata$_ZNKSt5ctypeIwE10do_toupperEPwPKw .text$_ZNKSt5ctypeIwE10do_tolowerEw .xdata$_ZNKSt5ctypeIwE10do_tolowerEw .pdata$_ZNKSt5ctypeIwE10do_tolowerEw .text$_ZNKSt5ctypeIwE10do_tolowerEPwPKw .xdata$_ZNKSt5ctypeIwE10do_tolowerEPwPKw .pdata$_ZNKSt5ctypeIwE10do_tolowerEPwPKw .text$_ZNKSt5ctypeIwE5do_isEtw .xdata$_ZNKSt5ctypeIwE5do_isEtw .pdata$_ZNKSt5ctypeIwE5do_isEtw .text$_ZNKSt5ctypeIwE5do_isEPKwS2_Pt .xdata$_ZNKSt5ctypeIwE5do_isEPKwS2_Pt .pdata$_ZNKSt5ctypeIwE5do_isEPKwS2_Pt .text$_ZNKSt5ctypeIwE10do_scan_isEtPKwS2_ .xdata$_ZNKSt5ctypeIwE10do_scan_isEtPKwS2_ .pdata$_ZNKSt5ctypeIwE10do_scan_isEtPKwS2_ .text$_ZNKSt5ctypeIwE11do_scan_notEtPKwS2_ .xdata$_ZNKSt5ctypeIwE11do_scan_notEtPKwS2_ .pdata$_ZNKSt5ctypeIwE11do_scan_notEtPKwS2_ .text$_ZNKSt5ctypeIwE8do_widenEc .xdata$_ZNKSt5ctypeIwE8do_widenEc .pdata$_ZNKSt5ctypeIwE8do_widenEc .text$_ZNKSt5ctypeIwE8do_widenEPKcS2_Pw .xdata$_ZNKSt5ct�      ypeIwE8do_widenEPKcS2_Pw .pdata$_ZNKSt5ctypeIwE8do_widenEPKcS2_Pw .text$_ZNKSt5ctypeIwE9do_narrowEwc .xdata$_ZNKSt5ctypeIwE9do_narrowEwc .pdata$_ZNKSt5ctypeIwE9do_narrowEwc .text$_ZNKSt5ctypeIwE9do_narrowEPKwS2_cPc .xdata$_ZNKSt5ctypeIwE9do_narrowEPKwS2_cPc .pdata$_ZNKSt5ctypeIwE9do_narrowEPKwS2_cPc .text$_ZNSt5ctypeIwE19_M_initialize_ctypeEv .xdata$_ZNSt5ctypeIwE19_M_initialize_ctypeEv .pdata$_ZNSt5ctypeIwE19_M_initialize_ctypeEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_decimal_pointEv _ZNKSt7__cxx1110moneypunctIcLb0EE16do_decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_thousands_sepEv _ZNKSt7__cxx1110moneypunctIcLb0EE16do_thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_frac_digitsEv _ZNKSt7__cxx1110moneypunctIcLb0EE14do_frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_pos_formatEv _ZNKSt7__cxx1110moneypunctIcLb0EE13do_pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_neg_formatEv _ZNKSt7__cxx1110moneypunctIcLb0EE13do_neg_formatEv .text$_ZNKSt7__cxx1110money�      punctIcLb1EE16do_decimal_pointEv _ZNKSt7__cxx1110moneypunctIcLb1EE16do_decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_thousands_sepEv _ZNKSt7__cxx1110moneypunctIcLb1EE16do_thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_frac_digitsEv _ZNKSt7__cxx1110moneypunctIcLb1EE14do_frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_pos_formatEv _ZNKSt7__cxx1110moneypunctIcLb1EE13do_pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_neg_formatEv _ZNKSt7__cxx1110moneypunctIcLb1EE13do_neg_formatEv .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED1Ev _ZNSt7__cxx1117moneypunct_bynameIcLb0EED1Ev .rdata$_ZTVNSt7__cxx1117moneypunct_bynameIcLb0EEE .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED1Ev _ZNSt7__cxx1117moneypunct_bynameIcLb1EED1Ev .rdata$_ZTVNSt7__cxx1117moneypunct_bynameIcLb1EEE .text$_ZNKSt7__cxx118numpunctIcE16do_decimal_pointEv _ZNKSt7__cxx118numpunctIcE16do_decimal_pointEv .text$_ZNKSt7__cxx118numpunctIcE16do_thousands_sepEv _ZNKSt7__cxx118numpunctIcE16do_thousands_sepEv .�      text$_ZNSt7__cxx1115numpunct_bynameIcED1Ev _ZNSt7__cxx1115numpunct_bynameIcED1Ev .rdata$_ZTVNSt7__cxx1115numpunct_bynameIcEE .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .text$_ZNKSt7__cxx118messagesIcE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale _ZNKSt7__cxx118messagesIcE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt7__cxx118messagesIcE8do_closeEi _ZNKSt7__cxx118messagesIcE8do_closeEi .text$_ZNKSt7__cxx117collateIcE7do_hashEPKcS3_ _ZNKSt7__cxx117collateIcE7do_hashEPKcS3_ .text$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7__cxx119money_putIcSt19�      ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED0Ev _ZNSt7__cxx1117moneypunct_bynameIcLb0EED0Ev .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED0Ev _ZNSt7__cxx1117moneypunct_bynameIcLb1EED0Ev .text$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_t�      raitsIcEEED0Ev .text$_ZNSt7__cxx1115numpunct_bynameIcED0Ev _ZNSt7__cxx1115numpunct_bynameIcED0Ev .text$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt7__cxx118messagesIcED1Ev _ZNSt7__cxx118messagesIcED1Ev .rdata$_ZTVNSt7__cxx118messagesIcEE .text$_ZNSt7__cxx118messagesIcED0Ev _ZNSt7__cxx118messagesIcED0Ev .text$_ZNSt7__cxx117collateIcED1Ev _ZNSt7__cxx117collateIcED1Ev .rdata$_ZTVNSt7__cxx117collateIcEE .text$_ZNSt7__cxx117collateIcED0Ev _ZNSt7__cxx117collateIcED0Ev .text$_ZNSt7__cxx1115messages_bynameIcED1Ev _ZNSt7__cxx1115messages_bynameIcED1Ev .text$_ZNSt7__cxx1115messages_bynameIcED0Ev _ZNSt7__cxx1115messages_bynameIcED0Ev .text$_ZNSt7__cxx1114collate_bynameIcED1Ev _ZNSt7__cxx1114collate_bynameIcED1Ev .text$_ZNSt7__cxx111�      4collate_bynameIcED0Ev _ZNSt7__cxx1114collate_bynameIcED0Ev .text$_ZNKSt7__cxx117collateIcE10do_compareEPKcS3_S3_S3_ _ZNKSt7__cxx117collateIcE10do_compareEPKcS3_S3_S3_ _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv.isra.33 .text$_ZNKSt7__cxx1110moneypunctIcLb1EE11do_groupingEv _ZNKSt7__cxx1110moneypunctIcLb1EE11do_groupingEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_curr_symbolEv _ZNKSt7__cxx1110moneypunctIcLb1EE14do_curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_positive_signEv _ZNKSt7__cxx1110moneypunctIcLb1EE16do_positive_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_negative_signEv _ZNKSt7__cxx1110moneypunctIcLb1EE16do_negative_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_curr_symbolEv _ZNKSt7__cxx1110moneypunctIcLb0EE14do_curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_positive_signEv _ZNKSt7__cxx1110moneypunctIcLb0EE16do_positive_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE11do_groupingEv _ZNKSt7__cxx1110moneypunctIcLb0EE11do_groupingEv .text$_ZNKSt�      7__cxx1110moneypunctIcLb0EE16do_negative_signEv _ZNKSt7__cxx1110moneypunctIcLb0EE16do_negative_signEv .text$_ZNKSt7__cxx118numpunctIcE11do_groupingEv _ZNKSt7__cxx118numpunctIcE11do_groupingEv .text$_ZNKSt7__cxx118numpunctIcE11do_truenameEv _ZNKSt7__cxx118numpunctIcE11do_truenameEv .text$_ZNKSt7__cxx118numpunctIcE12do_falsenameEv _ZNKSt7__cxx118numpunctIcE12do_falsenameEv .text$_ZNKSt7__cxx117collateIcE12do_transformEPKcS3_ _ZNKSt7__cxx117collateIcE12do_transformEPKcS3_ .text$_ZSt16__convert_from_vRKPiPciPKcz _ZSt16__convert_from_vRKPiPciPKcz .text$_ZNKSt5ctypeIcE5widenEPKcS2_Pc _ZNKSt5ctypeIcE5widenEPKcS2_Pc .text$_ZNSt7__cxx1110moneypunctIcLb0EEC2Ey _ZNSt7__cxx1110moneypunctIcLb0EEC2Ey .rdata$_ZTVNSt7__cxx1110moneypunctIcLb0EEE .text$_ZNSt7__cxx1110moneypunctIcLb0EEC1Ey _ZNSt7__cxx1110moneypunctIcLb0EEC1Ey .text$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy _ZNSt7__cxx1110moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .text$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPSt18__moneypunc�      t_cacheIcLb0EEy _ZNSt7__cxx1110moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .text$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPiPKcy _ZNSt7__cxx1110moneypunctIcLb0EEC2EPiPKcy .text$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPiPKcy _ZNSt7__cxx1110moneypunctIcLb0EEC1EPiPKcy .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13decimal_pointEv _ZNKSt7__cxx1110moneypunctIcLb0EE13decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13thousands_sepEv _ZNKSt7__cxx1110moneypunctIcLb0EE13thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE8groupingEv _ZNKSt7__cxx1110moneypunctIcLb0EE8groupingEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE11curr_symbolEv _ZNKSt7__cxx1110moneypunctIcLb0EE11curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13positive_signEv _ZNKSt7__cxx1110moneypunctIcLb0EE13positive_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE13negative_signEv _ZNKSt7__cxx1110moneypunctIcLb0EE13negative_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE11frac_digitsEv _ZNKSt7__cxx1110moneypunctIcLb0EE11frac_digitsEv .text$_ZNKSt7__cx�      x1110moneypunctIcLb0EE10pos_formatEv _ZNKSt7__cxx1110moneypunctIcLb0EE10pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIcLb0EE10neg_formatEv _ZNKSt7__cxx1110moneypunctIcLb0EE10neg_formatEv .text$_ZNSt7__cxx1110moneypunctIcLb1EEC2Ey _ZNSt7__cxx1110moneypunctIcLb1EEC2Ey .rdata$_ZTVNSt7__cxx1110moneypunctIcLb1EEE .text$_ZNSt7__cxx1110moneypunctIcLb1EEC1Ey _ZNSt7__cxx1110moneypunctIcLb1EEC1Ey .text$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEy _ZNSt7__cxx1110moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEy .text$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy _ZNSt7__cxx1110moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .text$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPiPKcy _ZNSt7__cxx1110moneypunctIcLb1EEC2EPiPKcy .text$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPiPKcy _ZNSt7__cxx1110moneypunctIcLb1EEC1EPiPKcy .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13decimal_pointEv _ZNKSt7__cxx1110moneypunctIcLb1EE13decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13thousands_sepEv _�      ZNKSt7__cxx1110moneypunctIcLb1EE13thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE8groupingEv _ZNKSt7__cxx1110moneypunctIcLb1EE8groupingEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE11curr_symbolEv _ZNKSt7__cxx1110moneypunctIcLb1EE11curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13positive_signEv _ZNKSt7__cxx1110moneypunctIcLb1EE13positive_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE13negative_signEv _ZNKSt7__cxx1110moneypunctIcLb1EE13negative_signEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE11frac_digitsEv _ZNKSt7__cxx1110moneypunctIcLb1EE11frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE10pos_formatEv _ZNKSt7__cxx1110moneypunctIcLb1EE10pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIcLb1EE10neg_formatEv _ZNKSt7__cxx1110moneypunctIcLb1EE10neg_formatEv .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2EPKcy _ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1EPKcy _ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb�      0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED2Ev _ZNSt7__cxx1117moneypunct_bynameIcLb0EED2Ev .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2EPKcy _ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1EPKcy _ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx111�      7moneypunct_bynameIcLb1EED2Ev _ZNSt7__cxx1117moneypunct_bynameIcLb1EED2Ev .text$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .text$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7__cxx119money_g�      etIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basece _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basece .text$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .text$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNKSt7__cxx119money_putIcSt19ostrea�      mbuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .data$_ZNSt7__cxx1110moneypunctIcLb1EE2idE .text$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .data$_ZNSt7__cxx1110moneypunctIcLb0EE2idE .text$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basece _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basece .text$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIc�      EEE6do_putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .text$_ZNSt7__cxx118numpunctIcEC2Ey _ZNSt7__cxx118numpunctIcEC2Ey .rdata$_ZTVNSt7__cxx118numpunctIcEE .text$_ZNSt7__cxx118numpunctIcEC1Ey _ZNSt7__cxx118numpunctIcEC1Ey .text$_ZNSt7__cxx118numpunctIcEC2EPSt16__numpunct_cacheIcEy _ZNSt7__cxx118numpunctIcEC2EPSt16__numpunct_cacheIcEy .text$_ZNSt7__cxx118numpunctIcEC1EPSt16__numpunct_cacheIcEy _ZNSt7__cxx118numpunctIcEC1EPSt16__numpunct_cacheIcEy .text$_ZNSt7__cxx118numpunctIcEC2EPiy _ZNSt7__cxx118numpunctIcEC2EPiy .text$_ZNSt7__cxx118numpunctIcEC1EPiy _ZNSt7__cxx118numpunctIcEC1EPiy .text$_ZNKSt7__cxx118numpunctIcE13decimal_pointEv _ZNKSt7__cxx118numpunctIcE13decimal_pointEv .text$_ZNKSt7__cxx118numpunctIcE13thousands_sepEv _ZNKSt7__cxx118numpunctIcE13thousands_sepEv .text$_ZNKSt7__cxx118numpunctIcE8groupingEv _ZNKSt7__cxx118numpunctIcE8groupingEv .text$_ZNKSt7__cxx118numpunctIcE8truenameEv _ZNKSt7__cxx118numpunctIcE8truenameEv .text$_ZNKSt7__cxx118numpunctIcE9falsenameEv _ZNKSt7__cxx118numpunct�      IcE9falsenameEv .text$_ZNSt7__cxx1115numpunct_bynameIcEC2EPKcy _ZNSt7__cxx1115numpunct_bynameIcEC2EPKcy .text$_ZNSt7__cxx1115numpunct_bynameIcEC1EPKcy _ZNSt7__cxx1115numpunct_bynameIcEC1EPKcy .text$_ZNSt7__cxx1115numpunct_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115numpunct_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115numpunct_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115numpunct_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115numpunct_bynameIcED2Ev _ZNSt7__cxx1115numpunct_bynameIcED2Ev .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .rdata$.refptr._ZTVSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC�      1ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .text$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNK�      St7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_trai�      tsIcEEED2Ev .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEE�      E14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .rdata$_ZTVNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNS_12basic_stringIcS3_SaIcEEEy _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNS_12basic_stringIcS3_SaIcEEEy .text$_ZNSt7__cxx1115t�      ime_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNS_12basic_stringIcS3_SaIcEEEy _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNS_12basic_stringIcS3_SaIcEEEy .text$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt7__cxx118messagesIcEC2Ey _ZNSt7__cxx118messagesIcEC2Ey .text$_ZNSt7__cxx118messagesIcEC1Ey _ZNSt7__cxx118messagesIcEC1Ey .text$_ZNSt7__cxx118messagesIcEC2EPiPKcy _ZNSt7__cxx118messagesIcEC2EPiPKcy .text$_ZNSt7__cxx118messagesIcEC1EPiPKcy _ZNSt7__cxx118messagesIcEC1EPiPKcy .text$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale _ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc _ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_trait�      sIcESaIcEEERKSt6localePKc .text$_ZNKSt7__cxx118messagesIcE3getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE _ZNKSt7__cxx118messagesIcE3getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNKSt7__cxx118messagesIcE5closeEi _ZNKSt7__cxx118messagesIcE5closeEi .text$_ZNSt7__cxx118messagesIcED2Ev _ZNSt7__cxx118messagesIcED2Ev .text$_ZNKSt7__cxx118messagesIcE18_M_convert_to_charERKNS_12basic_stringIcSt11char_traitsIcESaIcEEE _ZNKSt7__cxx118messagesIcE18_M_convert_to_charERKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNKSt7__cxx118messagesIcE20_M_convert_from_charEPc _ZNKSt7__cxx118messagesIcE20_M_convert_from_charEPc .text$_ZNSt7__cxx1115messages_bynameIcEC2EPKcy _ZNSt7__cxx1115messages_bynameIcEC2EPKcy .rdata$_ZTVNSt7__cxx1115messages_bynameIcEE .text$_ZNSt7__cxx1115messages_bynameIcEC1EPKcy _ZNSt7__cxx1115messages_bynameIcEC1EPKcy .text$_ZNSt7__cxx1115messages_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115messages_bynameIcEC2ERKNS_12basic_stringIcSt11char_�      traitsIcESaIcEEEy .text$_ZNSt7__cxx1115messages_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115messages_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115messages_bynameIcED2Ev _ZNSt7__cxx1115messages_bynameIcED2Ev _ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt12ctype_bynameIcEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt14codecvt_bynameIcciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt14codecvt_bynameIcciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .rdata$.refptr._ZTVSt14codecvt_bynameIcciE .text$_ZNSt14codecvt_bynameIcciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt14codecvt_bynameIcciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx117collateIcEC2Ey _ZNSt7__cxx117collateIcEC2Ey .text$_ZNSt7__cxx117collateIcEC1Ey _ZNSt7__cxx117collateIcEC1Ey .text$_ZNSt7__cxx117collateIcEC2EPiy _ZNSt7__cxx117collat�      eIcEC2EPiy .text$_ZNSt7__cxx117collateIcEC1EPiy _ZNSt7__cxx117collateIcEC1EPiy .text$_ZNKSt7__cxx117collateIcE7compareEPKcS3_S3_S3_ _ZNKSt7__cxx117collateIcE7compareEPKcS3_S3_S3_ .text$_ZNKSt7__cxx117collateIcE9transformEPKcS3_ _ZNKSt7__cxx117collateIcE9transformEPKcS3_ .text$_ZNKSt7__cxx117collateIcE4hashEPKcS3_ _ZNKSt7__cxx117collateIcE4hashEPKcS3_ .text$_ZNSt7__cxx117collateIcED2Ev _ZNSt7__cxx117collateIcED2Ev .text$_ZNSt7__cxx1114collate_bynameIcEC2EPKcy _ZNSt7__cxx1114collate_bynameIcEC2EPKcy .rdata$_ZTVNSt7__cxx1114collate_bynameIcEE .text$_ZNSt7__cxx1114collate_bynameIcEC1EPKcy _ZNSt7__cxx1114collate_bynameIcEC1EPKcy .text$_ZNSt7__cxx1114collate_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1114collate_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1114collate_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1114collate_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1114collate_bynameIcED2�      Ev _ZNSt7__cxx1114collate_bynameIcED2Ev .text$_ZSt9use_facetINSt7__cxx117collateIcEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx117collateIcEEERKT_RKSt6locale .data$_ZNSt7__cxx117collateIcE2idE .rdata$_ZTINSt7__cxx117collateIcEE .text$_ZSt9use_facetINSt7__cxx118numpunctIcEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118numpunctIcEEERKT_RKSt6locale .data$_ZNSt7__cxx118numpunctIcE2idE .rdata$_ZTINSt7__cxx118numpunctIcEE .text$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb1EEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx1110moneypunctIcLb1EEEERKT_RKSt6locale .rdata$_ZTINSt7__cxx1110moneypunctIcLb1EEE .text$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb0EEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx1110moneypunctIcLb0EEEERKT_RKSt6locale .rdata$_ZTINSt7__cxx1110moneypunctIcLb0EEE .text$_ZSt9use_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .data$_ZNSt7__cxx119money_putIcSt19ostream�      buf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZSt9use_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .data$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZSt9use_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .data$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .text$_ZSt9use_facetINSt7__cxx118messagesIcEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118messagesIcEEERKT_RKSt6locale .data$_ZNSt7__cxx118messagesIcE2idE .rdata�      $_ZTINSt7__cxx118messagesIcEE .text$_ZSt9has_facetINSt7__cxx117collateIcEEEbRKSt6locale _ZSt9has_facetINSt7__cxx117collateIcEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118numpunctIcEEEbRKSt6locale _ZSt9has_facetINSt7__cxx118numpunctIcEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx1110moneypunctIcLb0EEEEbRKSt6locale _ZSt9has_facetINSt7__cxx1110moneypunctIcLb0EEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118m�      essagesIcEEEbRKSt6locale _ZSt9has_facetINSt7__cxx118messagesIcEEEbRKSt6locale .text$_ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale _ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale .text$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKc _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .rdata$.refptr._ZNSt17__timepunct_cacheIcE12_S_timezonesE .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do�      _get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt�      12_Ios_IostateP2tmPKcSD_ _ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSD_ .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_base�      RSt12_Ios_IostateRe .text$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE _ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf�      _iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .data$_ZGVNSt7__cxx111�      0moneypunctIcLb0EE2idE .data$_ZGVNSt7__cxx1110moneypunctIcLb1EE2idE .data$_ZGVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt7__cxx118numpunctIcE2idE .data$_ZGVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt7__cxx118messagesIcE2idE .data$_ZGVNSt7__cxx117collateIcE2idE .rdata$_ZTSSt9time_base .rdata$_ZTISt9time_base .rdata$_ZTSSt10money_base .rdata$_ZTISt10money_base .rdata$_ZTSSt13messages_base .rdata$_ZTISt13messages_base .rdata$_ZTSNSt7__cxx117collateIcEE .rdata$_ZTSNSt7__cxx1114collate_bynameIcEE .rdata$_ZTINSt7__cxx1114collate_bynameIcEE .rdata$_ZTSNSt7__cxx118numpunctIcEE .rdata$_ZTSNSt7__cxx1115numpunct_bynameIcEE .rdata$_ZTINSt7__cxx1115numpunct_bynameIcEE .rdata$_ZTSNSt7__cxx1110moneypunctIcLb1EEE .rdata$_ZTSNSt7__cxx1110moneypunctIcLb0EEE .rdata$_ZTSNSt7__cxx118messagesIcEE .rdata$_ZTSNSt7__cxx1117moneypunct_bynameIcLb0EEE .rdata$_ZTIN�      St7__cxx1117moneypunct_bynameIcLb0EEE .rdata$_ZTSNSt7__cxx1117moneypunct_bynameIcLb1EEE .rdata$_ZTINSt7__cxx1117moneypunct_bynameIcLb1EEE .rdata$_ZTSNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .rdata$_ZTSNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE .rdata$_ZTSNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .rdata$_ZTSNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .rdata$_ZTINSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .rdata$_ZTSNSt7__cxx1115messages_bynameIcEE .rdata$_ZTINSt7__cxx1115messages_bynameIcEE .rdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EE4intlE .rdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EE4intlE .rdata$_ZNSt7__cxx1110moneypunctIcLb1EE4intlE .rdata$_ZNSt7__cxx1110moneypunctIcLb0EE4intlE .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_thousan�      ds_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13do_neg_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13do_neg_formatEv .x�      data$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED1Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED1Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED1Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED1Ev .xdata$_ZNKSt7__cxx118numpunctIcE16do_decimal_pointEv .pdata$_ZNKSt7__cxx118numpunctIcE16do_decimal_pointEv .xdata$_ZNKSt7__cxx118numpunctIcE16do_thousands_sepEv .pdata$_ZNKSt7__cxx118numpunctIcE16do_thousands_sepEv .xdata$_ZNSt7__cxx1115numpunct_bynameIcED1Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIcED1Ev .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .xdata$_ZNKSt7__cxx118messagesIcE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pdata$_ZNKSt7__cxx118messagesIcE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt7__cxx118messagesIcE8do_closeEi .pdata$_ZNKSt7__cxx118messagesIcE8do_closeEi .xdata$_ZNKSt7__cxx117collat�      eIcE7do_hashEPKcS3_ .pdata$_ZNKSt7__cxx117collateIcE7do_hashEPKcS3_ .xdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED0Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED0Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED0Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED0Ev .xdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEE�      ED0Ev .pdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt7__cxx1115numpunct_bynameIcED0Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIcED0Ev .xdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt7__cxx118messagesIcED1Ev .pdata$_ZNSt7__cxx118messagesIcED1Ev .xdata$_ZNSt7__cxx118messagesIcED0Ev .pdata$_ZNSt7__cxx118messagesIcED0Ev .xdata$_ZNSt7__cxx117collateIcED1Ev .pdata$_ZNSt7__cxx117collateIcED1Ev .xdata$_ZNSt7__cxx117collateIcED0Ev .pdata$_ZNSt7__cxx117collateIcED0Ev .xdata$_ZNSt7__cxx1115messages_bynameIcED1�      Ev .pdata$_ZNSt7__cxx1115messages_bynameIcED1Ev .xdata$_ZNSt7__cxx1115messages_bynameIcED0Ev .pdata$_ZNSt7__cxx1115messages_bynameIcED0Ev .xdata$_ZNSt7__cxx1114collate_bynameIcED1Ev .pdata$_ZNSt7__cxx1114collate_bynameIcED1Ev .xdata$_ZNSt7__cxx1114collate_bynameIcED0Ev .pdata$_ZNSt7__cxx1114collate_bynameIcED0Ev .xdata$_ZNKSt7__cxx117collateIcE10do_compareEPKcS3_S3_S3_ .pdata$_ZNKSt7__cxx117collateIcE10do_compareEPKcS3_S3_S3_ .text$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv.isra.33 .xdata$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv.isra.33 .pdata$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv.isra.33 .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11do_groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11do_groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE14do_curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_positive_signEv .xdata$_ZNKSt7__�      cxx1110moneypunctIcLb1EE16do_negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE16do_negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE14do_curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_positive_signEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11do_groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11do_groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE16do_negative_signEv .xdata$_ZNKSt7__cxx118numpunctIcE11do_groupingEv .pdata$_ZNKSt7__cxx118numpunctIcE11do_groupingEv .xdata$_ZNKSt7__cxx118numpunctIcE11do_truenameEv .pdata$_ZNKSt7__cxx118numpunctIcE11do_truenameEv .xdata$_ZNKSt7__cxx118numpunctIcE12do_falsenameEv .pdata$_ZNKSt7__cxx118numpunctIcE12do_falsenameEv .xdata$_ZNKSt7__cxx117collateIcE12do_transformEPKcS3_ .pdata$_ZNKSt7__cxx117collateIcE12do_transformEPKcS3_ .xdata$_ZSt16__convert_from_vRKP�      iPciPKcz .pdata$_ZSt16__convert_from_vRKPiPciPKcz .xdata$_ZNKSt5ctypeIcE5widenEPKcS2_Pc .pdata$_ZNKSt5ctypeIcE5widenEPKcS2_Pc .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2Ey .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2Ey .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1Ey .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1Ey .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC2EPiPKcy .xdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIcLb0EEC1EPiPKcy .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13thousa�      nds_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE8groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE8groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13positive_signEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE13negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE11frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE10pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE10pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb0EE10neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb0EE10neg_formatEv .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2Ey .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2Ey .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1Ey .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1Ey .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPSt18__m�      oneypunct_cacheIcLb1EEy .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEy .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC2EPiPKcy .xdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIcLb1EEC1EPiPKcy .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE8groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE8groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13positive_signEv .xdata$_ZN�      KSt7__cxx1110moneypunctIcLb1EE13negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE13negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE11frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE10pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE10pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIcLb1EE10neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIcLb1EE10neg_formatEv .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EEC1ERKNS_12basic_stringIcS�      t11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED2Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb0EED2Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED2Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIcLb1EED2Ev .xdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt7__cxx�      119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2E�      y .xdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basece .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basece .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_trait�      sIcEEE9_M_insertILb1EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES4_S4_RSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basece .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basece .xdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES4_bRSt8ios_basecRKNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNSt7__cxx118numpunctIcEC2Ey .pdata$_ZNSt7__cxx118numpunctIcEC2Ey .xdata$_ZNSt7__cxx118numpunctIcEC1Ey .pdata$_ZNSt7__cxx118numpunctIcEC1Ey .xdata$_ZNSt7__cxx118n�      umpunctIcEC2EPSt16__numpunct_cacheIcEy .pdata$_ZNSt7__cxx118numpunctIcEC2EPSt16__numpunct_cacheIcEy .xdata$_ZNSt7__cxx118numpunctIcEC1EPSt16__numpunct_cacheIcEy .pdata$_ZNSt7__cxx118numpunctIcEC1EPSt16__numpunct_cacheIcEy .xdata$_ZNSt7__cxx118numpunctIcEC2EPiy .pdata$_ZNSt7__cxx118numpunctIcEC2EPiy .xdata$_ZNSt7__cxx118numpunctIcEC1EPiy .pdata$_ZNSt7__cxx118numpunctIcEC1EPiy .xdata$_ZNKSt7__cxx118numpunctIcE13decimal_pointEv .pdata$_ZNKSt7__cxx118numpunctIcE13decimal_pointEv .xdata$_ZNKSt7__cxx118numpunctIcE13thousands_sepEv .pdata$_ZNKSt7__cxx118numpunctIcE13thousands_sepEv .xdata$_ZNKSt7__cxx118numpunctIcE8groupingEv .pdata$_ZNKSt7__cxx118numpunctIcE8groupingEv .xdata$_ZNKSt7__cxx118numpunctIcE8truenameEv .pdata$_ZNKSt7__cxx118numpunctIcE8truenameEv .xdata$_ZNKSt7__cxx118numpunctIcE9falsenameEv .pdata$_ZNKSt7__cxx118numpunctIcE9falsenameEv .xdata$_ZNSt7__cxx1115numpunct_bynameIcEC2EPKcy .pdata$_ZNSt7__cxx1115numpunct_bynameIcEC2EPKcy .xdata$_ZNSt7__cxx1115numpunct_bynameIcEC1EPKcy .pdata$_ZNSt7__cxx�      1115numpunct_bynameIcEC1EPKcy .xdata$_ZNSt7__cxx1115numpunct_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115numpunct_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115numpunct_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115numpunct_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115numpunct_bynameIcED2Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIcED2Ev .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNSt7__cxx1112basic_stringIcS2_SaIcEEEy .xdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iterat�      orIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_itera�      torIcSt11char_traitsIcEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_I�      os_Iostate .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf�      _iteratorIcSt11char_traitsIcEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNS_12basic_stringIcS3_SaIcEEEy .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKNS_12basic_stringIcS3_SaIcEEEy .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKNS_12basic_stringIcS3_SaIcEEEy .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iterator�      IcSt11char_traitsIcEEEC1ERKNS_12basic_stringIcS3_SaIcEEEy .xdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt7__cxx118messagesIcEC2Ey .pdata$_ZNSt7__cxx118messagesIcEC2Ey .xdata$_ZNSt7__cxx118messagesIcEC1Ey .pdata$_ZNSt7__cxx118messagesIcEC1Ey .xdata$_ZNSt7__cxx118messagesIcEC2EPiPKcy .pdata$_ZNSt7__cxx118messagesIcEC2EPiPKcy .xdata$_ZNSt7__cxx118messagesIcEC1EPiPKcy .pdata$_ZNSt7__cxx118messagesIcEC1EPiPKcy .xdata$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pdata$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc .pdata$_ZNKSt7__cxx118messagesIcE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc .xdata$_ZNKSt7__cxx118messagesIcE3getEiiiRKNS_12basic_stringIcSt11char�      _traitsIcESaIcEEE .pdata$_ZNKSt7__cxx118messagesIcE3getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNKSt7__cxx118messagesIcE5closeEi .pdata$_ZNKSt7__cxx118messagesIcE5closeEi .xdata$_ZNSt7__cxx118messagesIcED2Ev .pdata$_ZNSt7__cxx118messagesIcED2Ev .xdata$_ZNKSt7__cxx118messagesIcE18_M_convert_to_charERKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNKSt7__cxx118messagesIcE18_M_convert_to_charERKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNKSt7__cxx118messagesIcE20_M_convert_from_charEPc .pdata$_ZNKSt7__cxx118messagesIcE20_M_convert_from_charEPc .xdata$_ZNSt7__cxx1115messages_bynameIcEC2EPKcy .pdata$_ZNSt7__cxx1115messages_bynameIcEC2EPKcy .xdata$_ZNSt7__cxx1115messages_bynameIcEC1EPKcy .pdata$_ZNSt7__cxx1115messages_bynameIcEC1EPKcy .xdata$_ZNSt7__cxx1115messages_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115messages_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115messages_bynameIcEC1ERKNS_12basic_st�      ringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115messages_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115messages_bynameIcED2Ev .pdata$_ZNSt7__cxx1115messages_bynameIcED2Ev .text$_ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt14codecvt_bynameIcciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt14codecvt_bynameIcciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt14codecvt_bynameIcciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt14codecvt_bynameIcciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx117collateIcEC2Ey .pdata$_ZNSt7__cxx117collateIcEC2Ey .xdata$_ZNSt7__cxx117collateIcEC1Ey .pdata$_ZNSt7__cxx117collateIcEC1Ey .xdata$_ZNSt7__cxx117collat�      eIcEC2EPiy .pdata$_ZNSt7__cxx117collateIcEC2EPiy .xdata$_ZNSt7__cxx117collateIcEC1EPiy .pdata$_ZNSt7__cxx117collateIcEC1EPiy .xdata$_ZNKSt7__cxx117collateIcE7compareEPKcS3_S3_S3_ .pdata$_ZNKSt7__cxx117collateIcE7compareEPKcS3_S3_S3_ .xdata$_ZNKSt7__cxx117collateIcE9transformEPKcS3_ .pdata$_ZNKSt7__cxx117collateIcE9transformEPKcS3_ .xdata$_ZNKSt7__cxx117collateIcE4hashEPKcS3_ .pdata$_ZNKSt7__cxx117collateIcE4hashEPKcS3_ .xdata$_ZNSt7__cxx117collateIcED2Ev .pdata$_ZNSt7__cxx117collateIcED2Ev .xdata$_ZNSt7__cxx1114collate_bynameIcEC2EPKcy .pdata$_ZNSt7__cxx1114collate_bynameIcEC2EPKcy .xdata$_ZNSt7__cxx1114collate_bynameIcEC1EPKcy .pdata$_ZNSt7__cxx1114collate_bynameIcEC1EPKcy .xdata$_ZNSt7__cxx1114collate_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1114collate_bynameIcEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1114collate_bynameIcEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1114collate_bynameIcEC1ERKNS_12basic_stringIc�      St11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1114collate_bynameIcED2Ev .pdata$_ZNSt7__cxx1114collate_bynameIcED2Ev .xdata$_ZSt9use_facetINSt7__cxx117collateIcEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx117collateIcEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx118numpunctIcEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx118numpunctIcEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb1EEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb1EEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb0EEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx1110moneypunctIcLb0EEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx119money_getIcSt       19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx118messagesIcEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx118messagesIcEEERKT_RKSt6locale .xdata$_ZSt9has_facetINSt7__cxx117collateIcEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx117collateIcEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118numpunctIcEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx118numpunctIcEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx1110moneypunctIcLb0EEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx1110moneypunctIcLb0EEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx11      9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118messagesIcEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx118messagesIcEEEbRKSt6locale .xdata$_ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale .xdata$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ .pdata$_ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES4_S4_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES4_S4_RiPP      KcyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt7__cxx118time_getIcSt19istreamb      uf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSD_ .pdata$_ZNKSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSD_ .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEE      S4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .pdata$_ZNKSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS3_SaIcEEE .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cx      x11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_      ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIcS5_SaIcEEE _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKNSt7__cxx1112basic_stringIcSt11char_tra      itsIcESaIcEEERKSt6locale _ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIwS5_SaIwEEE _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEE _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKNSt7__cxx1112basic_stringIcS5_SaIcEEE _ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKNSt7__cxx1112basic_stringIwS5_SaIwEEE .text$_ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E       _ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .text$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E _ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .text$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ _ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .text$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ _ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .text$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ _ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb1EEPKNSt6locale5fa	      cetERNS_12__any_stringEPKT_SB_ .text$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ _ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1E
      EEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE _ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .text$_ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ _ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .text$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ _ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .text$_ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y _ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .text$_ZNSt13      __facet_shims14__messages_getIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y _ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .text$_ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi _ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .text$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi _ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .text$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE _ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .text$_ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE _ZNSt13__facet_shims20__time_get_dateorderIwE      ENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .text$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc _ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .text$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc _ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .text$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE _ZNSt13__facet_shims11__money_getIcEESt19istreambuf_      iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE _ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE _ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .text$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8      ios_baseS2_ePKNS_12__any_stringE _ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE _ZNKSt6locale5facet11_M_sso_shimEPKNS_2idE .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIcS5_SaIcEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIcS5_SaIcEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIcE6do_getESt19istreambuf_iteratorIcSt11char_traitsIcEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIcS5_SaIcEEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKNSt7__cxx      1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIwS5_SaIwEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIwS5_SaIwEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_get_shimIwE6do_getESt19istreambuf_iteratorIwSt11char_traitsIwEES6_bRSt8ios_baseRSt12_Ios_IostateRNSt7__cxx1112basic_stringIwS5_SaIwEEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pd      ata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE7do_openERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIcE6do_getEiiiRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_113messages_shimIwE6do_getEiiiRKNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKNS      t7__cxx1112basic_stringIcS5_SaIcEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKNSt7__cxx1112basic_stringIcS5_SaIcEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIcE6do_putESt19ostreambuf_iteratorIcSt11char_traitsIcEEbRSt8ios_basecRKNSt7__cxx1112basic_stringIcS5_SaIcEEE .text$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKNSt7__cxx1112basic_stringIwS5_SaIwEEE .xdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKNSt7__cxx1112basic_stringIwS5_SaIwEEE .pdata$_ZNKSt13__facet_shims12_GLOBAL__N_114money_put_shimIwE6do_putESt19ostreambuf_iteratorIwSt11char_traitsIwEEbRSt8ios_basewRKNSt7__cxx1112basic_stringIwS5_SaIwEEE .xdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .pdata$_ZNSt13__fa      cet_shims21__numpunct_fill_cacheIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .xdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .pdata$_ZNSt13__facet_shims21__numpunct_fill_cacheIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt16__numpunct_cacheIT_E .xdata$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .pdata$_ZNSt13__facet_shims17__collate_compareIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .xdata$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .pdata$_ZNSt13__facet_shims17__collate_compareIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKT_S9_S9_S9_ .xdata$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .pdata$_ZNSt13__facet_shims19__collate_transformIcEEvSt17integral_constantI      bLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .xdata$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .pdata$_ZNSt13__facet_shims19__collate_transformIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEPKT_SB_ .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIcLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdat      a$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb1EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .pdata$_ZNSt13__facet_shims23__moneypunct_fill_cacheIwLb0EEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEPSt18__moneypunct_cacheIT_XT0_EE .xdata$_ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .pdata$_ZNSt13__facet_shims15__messages_openIcEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .xdata$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .pdata$_ZNSt13__facet_shims15__messages_openIwEEiSt17integral_constantIbLb1EEPKNSt6locale5facetEPKcyRKS3_ .xdata$_ZNSt13__facet_shims14__messages_getIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .pdata$_ZNSt13__facet_shims14__messages_getIcEEvSt1      7integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .xdata$_ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .pdata$_ZNSt13__facet_shims14__messages_getIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetERNS_12__any_stringEiiiPKT_y .xdata$_ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .pdata$_ZNSt13__facet_shims16__messages_closeIcEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .xdata$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .pdata$_ZNSt13__facet_shims16__messages_closeIwEEvSt17integral_constantIbLb1EEPKNSt6locale5facetEi .xdata$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .pdata$_ZNSt13__facet_shims20__time_get_dateorderIcEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .xdata$_ZNSt13__facet_shims20__time_get_dateorderIwE      ENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .pdata$_ZNSt13__facet_shims20__time_get_dateorderIwEENSt9time_base9dateorderESt17integral_constantIbLb1EEPKNSt6locale5facetE .xdata$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .pdata$_ZNSt13__facet_shims10__time_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .xdata$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .pdata$_ZNSt13__facet_shims10__time_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_RSt8ios_baseRSt12_Ios_IostateP2tmc .xdata$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_co      nstantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_getIcEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_getIwEESt19istreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_S5_bRSt8ios_baseRSt12_Ios_IostatePePNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_putIcEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_eP      KNS_12__any_stringE .xdata$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .pdata$_ZNSt13__facet_shims11__money_putIwEESt19ostreambuf_iteratorIT_St11char_traitsIS2_EESt17integral_constantIbLb1EEPKNSt6locale5facetES5_bRSt8ios_baseS2_ePKNS_12__any_stringE .text$_ZNKSt6locale5facet11_M_sso_shimEPKNS_2idE .xdata$_ZNKSt6locale5facet11_M_sso_shimEPKNS_2idE .pdata$_ZNKSt6locale5facet11_M_sso_shimEPKNS_2idE .text$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_decimal_pointEv _ZNKSt7__cxx1110moneypunctIwLb0EE16do_decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_thousands_sepEv _ZNKSt7__cxx1110moneypunctIwLb0EE16do_thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE14do_frac_digitsEv _ZNKSt7__cxx1110moneypunctIwLb0EE14do_frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13do_pos_formatEv _ZNKSt7__cxx1110moneypunctIwLb0EE13do_pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13do      _neg_formatEv _ZNKSt7__cxx1110moneypunctIwLb0EE13do_neg_formatEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_decimal_pointEv _ZNKSt7__cxx1110moneypunctIwLb1EE16do_decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_thousands_sepEv _ZNKSt7__cxx1110moneypunctIwLb1EE16do_thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE14do_frac_digitsEv _ZNKSt7__cxx1110moneypunctIwLb1EE14do_frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_pos_formatEv _ZNKSt7__cxx1110moneypunctIwLb1EE13do_pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_neg_formatEv _ZNKSt7__cxx1110moneypunctIwLb1EE13do_neg_formatEv .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED1Ev _ZNSt7__cxx1117moneypunct_bynameIwLb0EED1Ev .rdata$_ZTVNSt7__cxx1117moneypunct_bynameIwLb0EEE .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED1Ev _ZNSt7__cxx1117moneypunct_bynameIwLb1EED1Ev .rdata$_ZTVNSt7__cxx1117moneypunct_bynameIwLb1EEE .text$_ZNKSt7__cxx118numpunctIwE16do_decimal_pointEv _ZNKSt7__cxx118numpunctIwE16do_decimal_pointEv .text$_ZN      KSt7__cxx118numpunctIwE16do_thousands_sepEv _ZNKSt7__cxx118numpunctIwE16do_thousands_sepEv .text$_ZNSt7__cxx1115numpunct_bynameIwED1Ev _ZNSt7__cxx1115numpunct_bynameIwED1Ev .rdata$_ZTVNSt7__cxx1115numpunct_bynameIwEE .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .text$_ZNKSt7__cxx118messagesIwE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale _ZNKSt7__cxx118messagesIwE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt7__cxx118messagesIwE8do_closeEi _ZNKSt7__cxx118messagesIwE8do_closeEi .text$_ZNKSt7__cxx117collateIwE7do_hashEPKwS3_ _ZNKSt7__cxx117collateIwE7do_hashEPKwS3_ .text$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZNSt7__cxx1      19money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED0Ev _ZNSt7__cxx1117moneypunct_bynameIwLb0EED0Ev .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED0Ev _ZNSt7__cxx1117moneypunct_bynameIwLb1EED0Ev .text$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt7__cxx119money_putIwSt19ostreambuf_ite      ratorIwSt11char_traitsIwEEED0Ev _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt7__cxx1115numpunct_bynameIwED0Ev _ZNSt7__cxx1115numpunct_bynameIwED0Ev .text$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt7__cxx118messagesIwED1Ev _ZNSt7__cxx118messagesIwED1Ev .rdata$_ZTVNSt7__cxx118messagesIwEE .text$_ZNSt7__cxx118messagesIwED0Ev _ZNSt7__cxx118messagesIwED0Ev .text$_ZNSt7__cxx117collateIwED1Ev _ZNSt7__cxx117collateIwED1Ev .rdata$_ZTVNSt7__cxx117collateIwEE .text$_ZNSt7__cxx117collateIwED0Ev _ZNSt7__cxx117collateIwED0Ev .text$_ZNSt7__cxx1115messages_bynameIwED1Ev _ZNSt7__cxx1115messages_bynameIwED1Ev .text$_ZNSt7__cxx1115messages_bynameIwED0Ev _ZNSt7__cxx1115messages_bynameIwED0Ev .text$_Z      NSt7__cxx1114collate_bynameIwED1Ev _ZNSt7__cxx1114collate_bynameIwED1Ev .text$_ZNSt7__cxx1114collate_bynameIwED0Ev _ZNSt7__cxx1114collate_bynameIwED0Ev .text$_ZNKSt7__cxx117collateIwE10do_compareEPKwS3_S3_S3_ _ZNKSt7__cxx117collateIwE10do_compareEPKwS3_S3_S3_ _ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.48 .text$_ZNKSt7__cxx1110moneypunctIwLb1EE11do_groupingEv _ZNKSt7__cxx1110moneypunctIwLb1EE11do_groupingEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE11do_groupingEv _ZNKSt7__cxx1110moneypunctIwLb0EE11do_groupingEv .text$_ZNKSt7__cxx118numpunctIwE11do_groupingEv _ZNKSt7__cxx118numpunctIwE11do_groupingEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_negative_signEv _ZNKSt7__cxx1110moneypunctIwLb1EE16do_negative_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE14do_curr_symbolEv _ZNKSt7__cxx1110moneypunctIwLb1EE14do_curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_positive_signEv _ZNKSt7__cxx1110moneypunctIwLb1EE16do_positive_signEv .text$_ZNKSt7__cxx118numpunctIwE12do_falsenameEv _ZNKS      t7__cxx118numpunctIwE12do_falsenameEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE14do_curr_symbolEv _ZNKSt7__cxx1110moneypunctIwLb0EE14do_curr_symbolEv .text$_ZNKSt7__cxx118numpunctIwE11do_truenameEv _ZNKSt7__cxx118numpunctIwE11do_truenameEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_positive_signEv _ZNKSt7__cxx1110moneypunctIwLb0EE16do_positive_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_negative_signEv _ZNKSt7__cxx1110moneypunctIwLb0EE16do_negative_signEv .text$_ZNKSt7__cxx117collateIwE12do_transformEPKwS3_ _ZNKSt7__cxx117collateIwE12do_transformEPKwS3_ .text$_ZNSt7__cxx1110moneypunctIwLb0EEC2Ey _ZNSt7__cxx1110moneypunctIwLb0EEC2Ey .rdata$_ZTVNSt7__cxx1110moneypunctIwLb0EEE .text$_ZNSt7__cxx1110moneypunctIwLb0EEC1Ey _ZNSt7__cxx1110moneypunctIwLb0EEC1Ey .text$_ZNSt7__cxx1110moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy _ZNSt7__cxx1110moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .text$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy _ZNSt7__cxx1110moneypunctIwLb0EEC1      EPSt18__moneypunct_cacheIwLb0EEy .text$_ZNSt7__cxx1110moneypunctIwLb0EEC2EPiPKcy _ZNSt7__cxx1110moneypunctIwLb0EEC2EPiPKcy .text$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPiPKcy _ZNSt7__cxx1110moneypunctIwLb0EEC1EPiPKcy .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13decimal_pointEv _ZNKSt7__cxx1110moneypunctIwLb0EE13decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13thousands_sepEv _ZNKSt7__cxx1110moneypunctIwLb0EE13thousands_sepEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE8groupingEv _ZNKSt7__cxx1110moneypunctIwLb0EE8groupingEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE11curr_symbolEv _ZNKSt7__cxx1110moneypunctIwLb0EE11curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13positive_signEv _ZNKSt7__cxx1110moneypunctIwLb0EE13positive_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE13negative_signEv _ZNKSt7__cxx1110moneypunctIwLb0EE13negative_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE11frac_digitsEv _ZNKSt7__cxx1110moneypunctIwLb0EE11frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE10pos_formatEv _ZNKSt7__cxx1       110moneypunctIwLb0EE10pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIwLb0EE10neg_formatEv _ZNKSt7__cxx1110moneypunctIwLb0EE10neg_formatEv .text$_ZNSt7__cxx1110moneypunctIwLb1EEC2Ey _ZNSt7__cxx1110moneypunctIwLb1EEC2Ey .rdata$_ZTVNSt7__cxx1110moneypunctIwLb1EEE .text$_ZNSt7__cxx1110moneypunctIwLb1EEC1Ey _ZNSt7__cxx1110moneypunctIwLb1EEC1Ey .text$_ZNSt7__cxx1110moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy _ZNSt7__cxx1110moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .text$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy _ZNSt7__cxx1110moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .text$_ZNSt7__cxx1110moneypunctIwLb1EEC2EPiPKcy _ZNSt7__cxx1110moneypunctIwLb1EEC2EPiPKcy .text$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPiPKcy _ZNSt7__cxx1110moneypunctIwLb1EEC1EPiPKcy .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13decimal_pointEv _ZNKSt7__cxx1110moneypunctIwLb1EE13decimal_pointEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13thousands_sepEv _ZNKSt7__cxx1110moneypunctIwLb1EE13thousands_sepEv !      .text$_ZNKSt7__cxx1110moneypunctIwLb1EE8groupingEv _ZNKSt7__cxx1110moneypunctIwLb1EE8groupingEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE11curr_symbolEv _ZNKSt7__cxx1110moneypunctIwLb1EE11curr_symbolEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13positive_signEv _ZNKSt7__cxx1110moneypunctIwLb1EE13positive_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE13negative_signEv _ZNKSt7__cxx1110moneypunctIwLb1EE13negative_signEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE11frac_digitsEv _ZNKSt7__cxx1110moneypunctIwLb1EE11frac_digitsEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE10pos_formatEv _ZNKSt7__cxx1110moneypunctIwLb1EE10pos_formatEv .text$_ZNKSt7__cxx1110moneypunctIwLb1EE10neg_formatEv _ZNKSt7__cxx1110moneypunctIwLb1EE10neg_formatEv .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2EPKcy _ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1EPKcy _ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcE"      EEy _ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED2Ev _ZNSt7__cxx1117moneypunct_bynameIwLb0EED2Ev .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2EPKcy _ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1EPKcy _ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1EPKcy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED2Ev _ZNSt7__cxx1117money#      punct_bynameIwLb1EED2Ev .text$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .text$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED$      2Ev .text$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewe _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewe .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .text$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1E%      EES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .data$_ZNSt7__cxx1110moneypunctIwLb1EE2idE .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .data$_ZNSt7__cxx1110moneypunctIwLb0EE2idE .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewe _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewe .text$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewRKNS_12basic_stringIwS&      3_SaIwEEE .text$_ZNSt7__cxx118numpunctIwEC2Ey _ZNSt7__cxx118numpunctIwEC2Ey .rdata$_ZTVNSt7__cxx118numpunctIwEE .text$_ZNSt7__cxx118numpunctIwEC1Ey _ZNSt7__cxx118numpunctIwEC1Ey .text$_ZNSt7__cxx118numpunctIwEC2EPSt16__numpunct_cacheIwEy _ZNSt7__cxx118numpunctIwEC2EPSt16__numpunct_cacheIwEy .text$_ZNSt7__cxx118numpunctIwEC1EPSt16__numpunct_cacheIwEy _ZNSt7__cxx118numpunctIwEC1EPSt16__numpunct_cacheIwEy .text$_ZNSt7__cxx118numpunctIwEC2EPiy _ZNSt7__cxx118numpunctIwEC2EPiy .text$_ZNSt7__cxx118numpunctIwEC1EPiy _ZNSt7__cxx118numpunctIwEC1EPiy .text$_ZNKSt7__cxx118numpunctIwE13decimal_pointEv _ZNKSt7__cxx118numpunctIwE13decimal_pointEv .text$_ZNKSt7__cxx118numpunctIwE13thousands_sepEv _ZNKSt7__cxx118numpunctIwE13thousands_sepEv .text$_ZNKSt7__cxx118numpunctIwE8groupingEv _ZNKSt7__cxx118numpunctIwE8groupingEv .text$_ZNKSt7__cxx118numpunctIwE8truenameEv _ZNKSt7__cxx118numpunctIwE8truenameEv .text$_ZNKSt7__cxx118numpunctIwE9falsenameEv _ZNKSt7__cxx118numpunctIwE9falsenameEv .text$_ZNSt7__cxx1115numpunct_byna'      meIwEC2EPKcy _ZNSt7__cxx1115numpunct_bynameIwEC2EPKcy .text$_ZNSt7__cxx1115numpunct_bynameIwEC1EPKcy _ZNSt7__cxx1115numpunct_bynameIwEC1EPKcy .text$_ZNSt7__cxx1115numpunct_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115numpunct_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115numpunct_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115numpunct_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115numpunct_bynameIwED2Ev _ZNSt7__cxx1115numpunct_bynameIwED2Ev .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .rdata$.refptr._ZTVSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEE(      y _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .text$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_it)      eratorIwSt11char_traitsIwEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNKSt7__cxx118time_*      getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES4_S4_RSt8ios_baseRS+      t12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .rdata$_ZTVNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNS_12basic_stringIcS2_IcESaIcEEEy _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNS_12basic_stringIcS2_IcESaIcEEEy .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_i,      teratorIwSt11char_traitsIwEEEC1ERKNS_12basic_stringIcS2_IcESaIcEEEy _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNS_12basic_stringIcS2_IcESaIcEEEy .text$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt7__cxx118messagesIwEC2Ey _ZNSt7__cxx118messagesIwEC2Ey .text$_ZNSt7__cxx118messagesIwEC1Ey _ZNSt7__cxx118messagesIwEC1Ey .text$_ZNSt7__cxx118messagesIwEC2EPiPKcy _ZNSt7__cxx118messagesIwEC2EPiPKcy .text$_ZNSt7__cxx118messagesIwEC1EPiPKcy _ZNSt7__cxx118messagesIwEC1EPiPKcy .text$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale _ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .text$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc _ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc -      .text$_ZNKSt7__cxx118messagesIwE3getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE _ZNKSt7__cxx118messagesIwE3getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .text$_ZNKSt7__cxx118messagesIwE5closeEi _ZNKSt7__cxx118messagesIwE5closeEi .text$_ZNSt7__cxx118messagesIwED2Ev _ZNSt7__cxx118messagesIwED2Ev .text$_ZNKSt7__cxx118messagesIwE18_M_convert_to_charERKNS_12basic_stringIwSt11char_traitsIwESaIwEEE _ZNKSt7__cxx118messagesIwE18_M_convert_to_charERKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .text$_ZNKSt7__cxx118messagesIwE20_M_convert_from_charEPc _ZNKSt7__cxx118messagesIwE20_M_convert_from_charEPc .text$_ZNSt7__cxx1115messages_bynameIwEC2EPKcy _ZNSt7__cxx1115messages_bynameIwEC2EPKcy .rdata$_ZTVNSt7__cxx1115messages_bynameIwEE .text$_ZNSt7__cxx1115messages_bynameIwEC1EPKcy _ZNSt7__cxx1115messages_bynameIwEC1EPKcy .text$_ZNSt7__cxx1115messages_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115messages_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_Z.      NSt7__cxx1115messages_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1115messages_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1115messages_bynameIwED2Ev _ZNSt7__cxx1115messages_bynameIwED2Ev _ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt12ctype_bynameIwEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt14codecvt_bynameIwciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt14codecvt_bynameIwciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .rdata$.refptr._ZTVSt14codecvt_bynameIwciE .text$_ZNSt14codecvt_bynameIwciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt14codecvt_bynameIwciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx117collateIwEC2Ey _ZNSt7__cxx117collateIwEC2Ey .text$_ZNSt7__cxx117collateIwEC1Ey _ZNSt7__cxx117collateIwEC1Ey .text$_ZNSt7__cxx117collateIwEC2EPiy _ZNSt7__cxx117collateIwEC2EPiy .text$_ZNSt7__c/      xx117collateIwEC1EPiy _ZNSt7__cxx117collateIwEC1EPiy .text$_ZNKSt7__cxx117collateIwE7compareEPKwS3_S3_S3_ _ZNKSt7__cxx117collateIwE7compareEPKwS3_S3_S3_ .text$_ZNKSt7__cxx117collateIwE9transformEPKwS3_ _ZNKSt7__cxx117collateIwE9transformEPKwS3_ .text$_ZNKSt7__cxx117collateIwE4hashEPKwS3_ _ZNKSt7__cxx117collateIwE4hashEPKwS3_ .text$_ZNSt7__cxx117collateIwED2Ev _ZNSt7__cxx117collateIwED2Ev .text$_ZNSt7__cxx1114collate_bynameIwEC2EPKcy _ZNSt7__cxx1114collate_bynameIwEC2EPKcy .rdata$_ZTVNSt7__cxx1114collate_bynameIwEE .text$_ZNSt7__cxx1114collate_bynameIwEC1EPKcy _ZNSt7__cxx1114collate_bynameIwEC1EPKcy .text$_ZNSt7__cxx1114collate_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1114collate_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1114collate_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy _ZNSt7__cxx1114collate_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZNSt7__cxx1114collate_bynameIwED2Ev _ZNSt7__cxx1114collate_0      bynameIwED2Ev .text$_ZSt9use_facetINSt7__cxx117collateIwEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx117collateIwEEERKT_RKSt6locale .data$_ZNSt7__cxx117collateIwE2idE .rdata$_ZTINSt7__cxx117collateIwEE .text$_ZSt9use_facetINSt7__cxx118numpunctIwEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118numpunctIwEEERKT_RKSt6locale .data$_ZNSt7__cxx118numpunctIwE2idE .rdata$_ZTINSt7__cxx118numpunctIwEE .text$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb1EEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx1110moneypunctIwLb1EEEERKT_RKSt6locale .rdata$_ZTINSt7__cxx1110moneypunctIwLb1EEE .text$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb0EEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx1110moneypunctIwLb0EEEERKT_RKSt6locale .rdata$_ZTINSt7__cxx1110moneypunctIwLb0EEE .text$_ZSt9use_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .data$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_tra1      itsIwEEE2idE .rdata$_ZTINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZSt9use_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .data$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZSt9use_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .data$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .text$_ZSt9use_facetINSt7__cxx118messagesIwEEERKT_RKSt6locale _ZSt9use_facetINSt7__cxx118messagesIwEEERKT_RKSt6locale .data$_ZNSt7__cxx118messagesIwE2idE .rdata$_ZTINSt7__cxx118messagesI2      wEE .text$_ZSt9has_facetINSt7__cxx117collateIwEEEbRKSt6locale _ZSt9has_facetINSt7__cxx117collateIwEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118numpunctIwEEEbRKSt6locale _ZSt9has_facetINSt7__cxx118numpunctIwEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx1110moneypunctIwLb0EEEEbRKSt6locale _ZSt9has_facetINSt7__cxx1110moneypunctIwLb0EEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale _ZSt9has_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .text$_ZSt9has_facetINSt7__cxx118messagesIwEEEbRKSt6locale _3      ZSt9has_facetINSt7__cxx118messagesIwEEEbRKSt6locale .text$_ZNKSt11__use_cacheISt16__numpunct_cacheIwEEclERKSt6locale _ZNKSt11__use_cacheISt16__numpunct_cacheIwEEclERKSt6locale .text$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE5equalERKS2_ _ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE5equalERKS2_ .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKw _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKw .rdata$.refptr._ZNSt17__timepunct_cacheIwE12_S_timezonesE .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES4_S4_RSt8ios_ba4      seRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_I5      ostateRNS_12basic_stringIcS2_IcESaIcEEE _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE _ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt86      ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istrea7      mbuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSD_ _ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSD_ _GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .data$_ZGVNSt7__cxx1110moneypunctIwL8      b0EE2idE .data$_ZGVNSt7__cxx1110moneypunctIwLb1EE2idE .data$_ZGVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt7__cxx118numpunctIwE2idE .data$_ZGVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt7__cxx118messagesIwE2idE .data$_ZGVNSt7__cxx117collateIwE2idE .rdata$_ZTSNSt7__cxx117collateIwEE .rdata$_ZTSNSt7__cxx1114collate_bynameIwEE .rdata$_ZTINSt7__cxx1114collate_bynameIwEE .rdata$_ZTSNSt7__cxx118numpunctIwEE .rdata$_ZTSNSt7__cxx1115numpunct_bynameIwEE .rdata$_ZTINSt7__cxx1115numpunct_bynameIwEE .rdata$_ZTSNSt7__cxx1110moneypunctIwLb1EEE .rdata$_ZTSNSt7__cxx1110moneypunctIwLb0EEE .rdata$_ZTSNSt7__cxx118messagesIwEE .rdata$_ZTSNSt7__cxx1117moneypunct_bynameIwLb0EEE .rdata$_ZTINSt7__cxx1117moneypunct_bynameIwLb0EEE .rdata$_ZTSNSt7__cxx1117moneypunct_bynameIwLb1EEE .rdata$_ZTINSt7__cxx1117moneypunct_bynameIwLb1EEE .rdata$_ZTSNSt7__cxx119money_getIw9      St19istreambuf_iteratorIwSt11char_traitsIwEEEE .rdata$_ZTSNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE .rdata$_ZTSNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .rdata$_ZTSNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .rdata$_ZTINSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .rdata$_ZTSNSt7__cxx1115messages_bynameIwEE .rdata$_ZTINSt7__cxx1115messages_bynameIwEE .rdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EE4intlE .rdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EE4intlE .rdata$_ZNSt7__cxx1110moneypunctIwLb1EE4intlE .rdata$_ZNSt7__cxx1110moneypunctIwLb0EE4intlE .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE14do_frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE14d:      o_frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13do_pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13do_pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13do_neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13do_neg_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE14do_frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE14do_frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13do_neg_formatEv .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED1Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED1Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED1Ev .pdata$_ZNSt7__cxx111;      7moneypunct_bynameIwLb1EED1Ev .xdata$_ZNKSt7__cxx118numpunctIwE16do_decimal_pointEv .pdata$_ZNKSt7__cxx118numpunctIwE16do_decimal_pointEv .xdata$_ZNKSt7__cxx118numpunctIwE16do_thousands_sepEv .pdata$_ZNKSt7__cxx118numpunctIwE16do_thousands_sepEv .xdata$_ZNSt7__cxx1115numpunct_bynameIwED1Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIwED1Ev .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .xdata$_ZNKSt7__cxx118messagesIwE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pdata$_ZNKSt7__cxx118messagesIwE7do_openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt7__cxx118messagesIwE8do_closeEi .pdata$_ZNKSt7__cxx118messagesIwE8do_closeEi .xdata$_ZNKSt7__cxx117collateIwE7do_hashEPKwS3_ .pdata$_ZNKSt7__cxx117collateIwE7do_hashEPKwS3_ .xdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7__cxx119m<      oney_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED0Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED0Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED0Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED0Ev .xdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .p=      data$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt7__cxx1115numpunct_bynameIwED0Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIwED0Ev .xdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt7__cxx118messagesIwED1Ev .pdata$_ZNSt7__cxx118messagesIwED1Ev .xdata$_ZNSt7__cxx118messagesIwED0Ev .pdata$_ZNSt7__cxx118messagesIwED0Ev .xdata$_ZNSt7__cxx117collateIwED1Ev .pdata$_ZNSt7__cxx117collateIwED1Ev .xdata$_ZNSt7__cxx117collateIwED0Ev .pdata$_ZNSt7__cxx117collateIwED0Ev .xdata$_ZNSt7__cxx1115messages_bynameIwED1Ev .pdata$_ZNSt7__cxx1115messages_bynameIwED1Ev .xdata$_ZNSt7__cxx1115messages_bynameIwED0Ev .pdata$_ZNSt7__cxx1115messages_bynameIwED0Ev .xdata$_ZNSt7__cxx1114collate_byna>      meIwED1Ev .pdata$_ZNSt7__cxx1114collate_bynameIwED1Ev .xdata$_ZNSt7__cxx1114collate_bynameIwED0Ev .pdata$_ZNSt7__cxx1114collate_bynameIwED0Ev .xdata$_ZNKSt7__cxx117collateIwE10do_compareEPKwS3_S3_S3_ .pdata$_ZNKSt7__cxx117collateIwE10do_compareEPKwS3_S3_S3_ .text$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.48 .xdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.48 .pdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.48 .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11do_groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11do_groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11do_groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11do_groupingEv .xdata$_ZNKSt7__cxx118numpunctIwE11do_groupingEv .pdata$_ZNKSt7__cxx118numpunctIwE11do_groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE14do_curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb?      1EE14do_curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE16do_positive_signEv .xdata$_ZNKSt7__cxx118numpunctIwE12do_falsenameEv .pdata$_ZNKSt7__cxx118numpunctIwE12do_falsenameEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE14do_curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE14do_curr_symbolEv .xdata$_ZNKSt7__cxx118numpunctIwE11do_truenameEv .pdata$_ZNKSt7__cxx118numpunctIwE11do_truenameEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_positive_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE16do_negative_signEv .xdata$_ZNKSt7__cxx117collateIwE12do_transformEPKwS3_ .pdata$_ZNKSt7__cxx117collateIwE12do_transformEPKwS3_ .xdata$_ZNSt7__cxx1110moneypunctIwLb0EEC2Ey .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC2Ey .xdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1Ey .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1Ey .xdata$_ZNSt7__cxx1110moneyp@      unctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .xdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy .xdata$_ZNSt7__cxx1110moneypunctIwLb0EEC2EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC2EPiPKcy .xdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIwLb0EEC1EPiPKcy .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE8groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE8groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13posiA      tive_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE13negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE11frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE10pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE10pos_formatEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb0EE10neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb0EE10neg_formatEv .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC2Ey .pdata$_ZNSt7__cxx1110moneypunctIwLb1EEC2Ey .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1Ey .pdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1Ey .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .pdata$_ZNSt7__cxx1110moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .pdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC2EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIwLB      b1EEC2EPiPKcy .xdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPiPKcy .pdata$_ZNSt7__cxx1110moneypunctIwLb1EEC1EPiPKcy .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13decimal_pointEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13decimal_pointEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13thousands_sepEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13thousands_sepEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE8groupingEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE8groupingEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11curr_symbolEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11curr_symbolEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13positive_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13positive_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13negative_signEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE13negative_signEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11frac_digitsEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE11frac_digitsEv .xdata$_ZNKSt7__cxx1110moneypunctIwLb1EE10pos_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE10pos_formatEv .xC      data$_ZNKSt7__cxx1110moneypunctIwLb1EE10neg_formatEv .pdata$_ZNKSt7__cxx1110moneypunctIwLb1EE10neg_formatEv .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED2Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb0EED2Ev .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1EPKcy .pdata$_ZNSt7__cxx1117moneypunct_bynameID      wLb1EEC1EPKcy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED2Ev .pdata$_ZNSt7__cxx1117moneypunct_bynameIwLb1EED2Ev .xdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11E      char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewe .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11F      char_traitsIwEEE3putES4_bRSt8ios_basewe .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES4_S4_RSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES4_S4_RSt8ios_bG      asewRKNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewe .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewe .xdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES4_bRSt8ios_basewRKNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNSt7__cxx118numpunctIwEC2Ey .pdata$_ZNSt7__cxx118numpunctIwEC2Ey .xdata$_ZNSt7__cxx118numpunctIwEC1Ey .pdata$_ZNSt7__cxx118numpunctIwEC1Ey .xdata$_ZNSt7__cxx118numpunctIwEC2EPSt16__numpunct_cacheIwEy .pdata$_ZNSt7__cxx118numpunctIwEC2EPSt16__numpunct_cacheIwEy .xdata$_ZNSt7__cxx118numpunctIwEC1EPSt16__numpunct_cacheIwEy .pdata$_ZNSt7__cxx118numpunctIwEC1EPSt16__numpunct_cacheIwEy .xdata$_ZNSt7__cxx118numpunctIwEC2EPiy .pdata$_ZNSt7__cxx118numpunctIwEC2EPiy .xdata$_ZNSt7__cxx118numpunctIH      wEC1EPiy .pdata$_ZNSt7__cxx118numpunctIwEC1EPiy .xdata$_ZNKSt7__cxx118numpunctIwE13decimal_pointEv .pdata$_ZNKSt7__cxx118numpunctIwE13decimal_pointEv .xdata$_ZNKSt7__cxx118numpunctIwE13thousands_sepEv .pdata$_ZNKSt7__cxx118numpunctIwE13thousands_sepEv .xdata$_ZNKSt7__cxx118numpunctIwE8groupingEv .pdata$_ZNKSt7__cxx118numpunctIwE8groupingEv .xdata$_ZNKSt7__cxx118numpunctIwE8truenameEv .pdata$_ZNKSt7__cxx118numpunctIwE8truenameEv .xdata$_ZNKSt7__cxx118numpunctIwE9falsenameEv .pdata$_ZNKSt7__cxx118numpunctIwE9falsenameEv .xdata$_ZNSt7__cxx1115numpunct_bynameIwEC2EPKcy .pdata$_ZNSt7__cxx1115numpunct_bynameIwEC2EPKcy .xdata$_ZNSt7__cxx1115numpunct_bynameIwEC1EPKcy .pdata$_ZNSt7__cxx1115numpunct_bynameIwEC1EPKcy .xdata$_ZNSt7__cxx1115numpunct_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115numpunct_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115numpunct_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115numpuI      nct_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115numpunct_bynameIwED2Ev .pdata$_ZNSt7__cxx1115numpunct_bynameIwED2Ev .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNSt7__cxx1112basic_stringIcS1_IcESaIcEEEy .xdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt7__cxx118time_getIwSt19istreambufJ      _iteratorIwSt11char_traitsIwEEE10date_orderEv .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES4_S4_RSt8ios_bK      aseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES4_S4_RiiiyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreL      ambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy M      .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNS_12basic_stringIcS2_IcESaIcEEEy .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKNS_12basic_stringIcS2_IcESaIcEEEy .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNS_12basic_stringIcS2_IcESaIcEEEy .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKNS_12basic_stringIcS2_IcESaIcEEEy .xdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt7__cxx118messagesIwEC2Ey .pdata$_ZNSt7__cxx118messagesIwECN      2Ey .xdata$_ZNSt7__cxx118messagesIwEC1Ey .pdata$_ZNSt7__cxx118messagesIwEC1Ey .xdata$_ZNSt7__cxx118messagesIwEC2EPiPKcy .pdata$_ZNSt7__cxx118messagesIwEC2EPiPKcy .xdata$_ZNSt7__cxx118messagesIwEC1EPiPKcy .pdata$_ZNSt7__cxx118messagesIwEC1EPiPKcy .xdata$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .pdata$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6locale .xdata$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc .pdata$_ZNKSt7__cxx118messagesIwE4openERKNS_12basic_stringIcSt11char_traitsIcESaIcEEERKSt6localePKc .xdata$_ZNKSt7__cxx118messagesIwE3getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .pdata$_ZNKSt7__cxx118messagesIwE3getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .xdata$_ZNKSt7__cxx118messagesIwE5closeEi .pdata$_ZNKSt7__cxx118messagesIwE5closeEi .xdata$_ZNSt7__cxx118messagesIwED2Ev .pdata$_ZNSt7__cxx118messagesIwED2Ev .xdata$_ZNKSt7__cxx118messagesIwE18_M_convO      ert_to_charERKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .pdata$_ZNKSt7__cxx118messagesIwE18_M_convert_to_charERKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .xdata$_ZNKSt7__cxx118messagesIwE20_M_convert_from_charEPc .pdata$_ZNKSt7__cxx118messagesIwE20_M_convert_from_charEPc .xdata$_ZNSt7__cxx1115messages_bynameIwEC2EPKcy .pdata$_ZNSt7__cxx1115messages_bynameIwEC2EPKcy .xdata$_ZNSt7__cxx1115messages_bynameIwEC1EPKcy .pdata$_ZNSt7__cxx1115messages_bynameIwEC1EPKcy .xdata$_ZNSt7__cxx1115messages_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115messages_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115messages_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1115messages_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1115messages_bynameIwED2Ev .pdata$_ZNSt7__cxx1115messages_bynameIwED2Ev .text$_ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdatP      a$_ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt14codecvt_bynameIwciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt14codecvt_bynameIwciEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt14codecvt_bynameIwciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt14codecvt_bynameIwciEC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx117collateIwEC2Ey .pdata$_ZNSt7__cxx117collateIwEC2Ey .xdata$_ZNSt7__cxx117collateIwEC1Ey .pdata$_ZNSt7__cxx117collateIwEC1Ey .xdata$_ZNSt7__cxx117collateIwEC2EPiy .pdata$_ZNSt7__cxx117collateIwEC2EPiy .xdata$_ZNSt7__cxx117collateIwEC1EPiy .pdata$_ZNSt7__cxx117collateIwEC1EPiy .xdata$_ZNKSt7__cxx117collateIwE7compareEPKwS3_S3_S3_ .pdata$_ZNKSt7__cxx117collateIwE7compareEPKwS3_S3_S3_ .xdata$_ZNKSt7__cxx117collateIwE9transformEPKwS3_ .pdata$_ZNKSt7__cxx117cQ      ollateIwE9transformEPKwS3_ .xdata$_ZNKSt7__cxx117collateIwE4hashEPKwS3_ .pdata$_ZNKSt7__cxx117collateIwE4hashEPKwS3_ .xdata$_ZNSt7__cxx117collateIwED2Ev .pdata$_ZNSt7__cxx117collateIwED2Ev .xdata$_ZNSt7__cxx1114collate_bynameIwEC2EPKcy .pdata$_ZNSt7__cxx1114collate_bynameIwEC2EPKcy .xdata$_ZNSt7__cxx1114collate_bynameIwEC1EPKcy .pdata$_ZNSt7__cxx1114collate_bynameIwEC1EPKcy .xdata$_ZNSt7__cxx1114collate_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1114collate_bynameIwEC2ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1114collate_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .pdata$_ZNSt7__cxx1114collate_bynameIwEC1ERKNS_12basic_stringIcSt11char_traitsIcESaIcEEEy .xdata$_ZNSt7__cxx1114collate_bynameIwED2Ev .pdata$_ZNSt7__cxx1114collate_bynameIwED2Ev .xdata$_ZSt9use_facetINSt7__cxx117collateIwEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx117collateIwEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx118numpunctIwEEERKT_RKSt6locale .pdaR      ta$_ZSt9use_facetINSt7__cxx118numpunctIwEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb1EEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb1EEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb0EEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx1110moneypunctIwLb0EEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEERKT_RKSt6locale .xdata$_ZSt9use_facetINSt7__cxxS      118messagesIwEEERKT_RKSt6locale .pdata$_ZSt9use_facetINSt7__cxx118messagesIwEEERKT_RKSt6locale .xdata$_ZSt9has_facetINSt7__cxx117collateIwEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx117collateIwEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118numpunctIwEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx118numpunctIwEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx1110moneypunctIwLb0EEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx1110moneypunctIwLb0EEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .pdata$_ZSt9has_facetINStT      7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEEbRKSt6locale .xdata$_ZSt9has_facetINSt7__cxx118messagesIwEEEbRKSt6locale .pdata$_ZSt9has_facetINSt7__cxx118messagesIwEEEbRKSt6locale .xdata$_ZNKSt11__use_cacheISt16__numpunct_cacheIwEEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt16__numpunct_cacheIwEEclERKSt6locale .xdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE5equalERKS2_ .pdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE5equalERKS2_ .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES4_S4_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKw .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES4_S4_RSt8ios_baseRSt12_Ios_U      IostateP2tmPKw .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_basV      eRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES4_S4_S4_RSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIcS2_IcESaIcEEE .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11chaW      r_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .pdata$_ZNKSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES4_S4_bRSt8ios_baseRSt12_Ios_IostateRNS_12basic_stringIwS3_SaIwEEE .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx1X      1IjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11ImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intB5cxx11IyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSD_ .pdata$_ZNKSt7__cxxY      118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES4_S4_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSD_ .text.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .xdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .pdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEy .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED1Ev _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED1Ev .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED1Ev _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED1Ev .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED0Ev _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED0Ev .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv _ZN9__gnu_Z      cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4syncEv _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4syncEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_Seek[      dirSt13_Ios_Openmode _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE5uflowEv _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE5uflowEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsgetnEPwx _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsgetnEPwx .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9underflowEv _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9underflowEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9pbackfailEt _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9pbackfailEt .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE8overflowEt _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE8overflowEt .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsputnEPKwx _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsputnEPKwx .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsputnEP\      Kcx _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsputnEPKcx .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcx _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcx .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED1Ev _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED1Ev .rdata$.refptr._ZTVSt13basic_filebufIwSt11char_traitsIwEE .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED1Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED1Ev .rdata$.refptr._ZTVSt13basic_filebufIcSt11char_traitsIcEE .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED0Ev _ZN9__gnu_cxx13stdio_filebu]      fIcSt11char_traitsIcEED0Ev .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED0Ev _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED0Ev .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev .rdata$_ZTVN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1Ev .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EiSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EiSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP6_iobufSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP6_iobufSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EP6_iobufSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIcSt11char^      _traitsIcEEC1EP6_iobufSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4swapERS3_ _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4swapERS3_ .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv .text$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP6_iobuf _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP6_iobuf .rdata$_ZTVN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EP6_iobuf _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EP6_iobuf .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EOS3_ .text$_ZN9__gnu_cxx18stdio_s_      ync_filebufIcSt11char_traitsIcEEC1EOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EOS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEaSEOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEaSEOS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4swapERS3_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4swapERS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2Ev _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2Ev .rdata$_ZTVN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1Ev _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1Ev .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EiSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EiSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EiSt13_Ios_Openmodey _Z`      N9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EiSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EP6_iobufSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EP6_iobufSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EP6_iobufSt13_Ios_Openmodey _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EP6_iobufSt13_Ios_Openmodey .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED2Ev _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED2Ev .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4swapERS3_ _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4swapERS3_ .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE2fdEv _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE2fdEv .text$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4fileEv _ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4fileEv .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EP6_iobuf _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EP6_iobuf .rdaa      ta$_ZTVN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EP6_iobuf _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EP6_iobuf .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EOS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EOS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEaSEOS3_ _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEaSEOS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4swapERS3_ _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4swapERS3_ .text$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4fileEv _ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4fileEv .rdata$_ZTSN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE .rdata$_ZTIN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE .rdata$_ZTSN9__gnu_cxx18stdio_sb      ync_filebufIwSt11char_traitsIwEEE .rdata$_ZTIN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE .rdata$_ZTSN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE .rdata$_ZTIN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE .rdata$_ZTSN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE .rdata$_ZTIN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED1Ev .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED1Ev .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED1Ev .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED1Ev .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED0Ev .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEED0Ev .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv .xdata$_Zc      N9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4syncEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4syncEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Od      penmode .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE5uflowEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE5uflowEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsgetnEPwx .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsgetnEPwx .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9underflowEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9underflowEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9pbackfailEt .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE9pbackfailEt .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE8overflowEt .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE8overflowEt .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsputnEPKwx .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE6xsputnEPKwx .xdata$_ZN9__gnu_cxx18stdioe      _sync_filebufIcSt11char_traitsIcEE6xsputnEPKcx .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsputnEPKcx .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcx .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcx .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED1Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED1Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED1Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED1Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED0Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsf      IcEED0Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED0Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED0Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EiSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EiSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP6_iobufSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP6_iobufSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EP6_iobufSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EP6_iobufg      St13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4swapERS3_ .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4swapERS3_ .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv .xdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv .pdata$_ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP6_iobuf .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP6_iobuf .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EP6_iobuf .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EP6_iobuf .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIch      EEC1EOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEaSEOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEaSEOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4swapERS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4swapERS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EiSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EiSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EiSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIi      wSt11char_traitsIwEEC1EiSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EP6_iobufSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC2EP6_iobufSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EP6_iobufSt13_Ios_Openmodey .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEC1EP6_iobufSt13_Ios_Openmodey .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED2Ev .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEED2Ev .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4swapERS3_ .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4swapERS3_ .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE2fdEv .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE2fdEv .xdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4fileEv .pdata$_ZN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEE4fileEv .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EP6_iobuf .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11chj      ar_traitsIwEEC2EP6_iobuf .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EP6_iobuf .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EP6_iobuf .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC2EOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEC1EOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEaSEOS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEaSEOS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4swapERS3_ .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4swapERS3_ .xdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4fileEv .pdata$_ZN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEE4fileEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcx _ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcx .text$_ZNSt13basic_filebufIwSt11char_k      traitsIwEE6setbufEPwx _ZNSt13basic_filebufIwSt11char_traitsIwEE6setbufEPwx .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv _ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE9showmanycEv _ZNSt13basic_filebufIwSt11char_traitsIwEE9showmanycEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv _ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE4syncEv _ZNSt13basic_filebufIwSt11char_traitsIwEE4syncEv _ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv.part.41 .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi _ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE9pbackfailEt _ZNSt13basic_filebufIwSt11char_traitsIwEE9pbackfailEt .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv _ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE9underflowEv _ZNSt13basic_filebufIwl      St11char_traitsIwEE9underflowEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcx _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcx .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsputnEPKwx _ZNSt13basic_filebufIwSt11char_traitsIwEE6xsputnEPKwx .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcx _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcx .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsgetnEPwx _ZNSt13basic_filebufIwSt11char_traitsIwEE6xsgetnEPwx .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv _ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv _ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev _ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev .rdata$_ZTVSt13basic_filebufIcSt11char_traitsIcEE .text$_ZNSt13basic_filebufIcSt11char_traitsIcEEC1Ev _ZNSt13basic_filebufIcSt11char_traitsIcEEC1Ev .text$_ZNSt13basic_filebufIcm      St11char_traitsIcEEC2EOS2_ _ZNSt13basic_filebufIcSt11char_traitsIcEEC2EOS2_ .text$_ZNSt13basic_filebufIcSt11char_traitsIcEEC1EOS2_ _ZNSt13basic_filebufIcSt11char_traitsIcEEC1EOS2_ .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE4swapERS2_ _ZNSt13basic_filebufIcSt11char_traitsIcEE4swapERS2_ .text$_ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv _ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv _ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv _ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcx _ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcx .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posERi _ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posERi .text$_ZNSt13basic_filebufIcSt11char_tn      raitsIcEE19_M_terminate_outputEv _ZNSt13basic_filebufIcSt11char_traitsIcEE19_M_terminate_outputEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdiri _ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdiri .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi _ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE13_M_set_bufferEx _ZNSt13basic_filebufIcSt11char_traitsIcEE13_M_set_bufferEx .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EOS2_ _ZNSt14basic_ifstro      eamIcSt11char_traitsIcEEC2EOS2_ .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EOS2_ _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EOS2_ .rdata$_ZTCSt14basic_ifstreamIcSt11char_traitsIcEE0_Si .rdata$_ZTVSt14basic_ifstreamIcSt11char_traitsIcEE .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4swapERS2_ _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4swapERS2_ .text$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv _ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EOS2_ _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EOS2_ .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EOS2_ _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EOS2_ .rdata$_ZTCSt14basic_ofstreamIcSt11char_traitsIcEE0_So .rdata$_ZTVSt14basic_ofstreamIcSt11char_traitsIcEE .text$p      _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4swapERS2_ _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4swapERS2_ .text$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EOS2_ _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EOS2_ .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EOS2_ _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EOS2_ .rdata$_ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Si .rdata$_ZTVSt13basic_fstreamIcSt11char_traitsIcEE .rdata$_ZTCSt13basic_fstreamIcSt11char_traitsIcEE16_So .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4swapERS2_ _ZNSt13basic_fstreamIcSt11char_traitsIcEE4swapERS2_ .text$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE5rdbufEv _ZNKSt13basic_fstreamIcSt11char_traitsIcq      EE5rdbufEv .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _ZNSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE15_M_create_pbackEv _ZNSt13basic_filebufIwSt11char_traitsIwEE15_M_create_pbackEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE16_M_destroy_pbackEv _ZNSt13basic_filebufIwSt11char_traitsIwEE16_M_destroy_pbackEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2Ev _ZNSt13basic_filebufIwSt11char_traitsIwEEC2Ev .rdata$_ZTVSt13basic_filebufIwSt11char_traitsIwEE .text$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1Ev _ZNSt13basic_filebufIwSt11char_traitsIwEEC1Ev .text$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2EOS2_ _ZNSt13basic_filebufIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1EOS2_ _ZNSt13basic_filebufIwSt11char_traitsIwEEC1EOS2_ .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE4swapERS2_ _ZNSt13basic_r      filebufIwSt11char_traitsIwEE4swapERS2_ .text$_ZNKSt13basic_filebufIwSt11char_traitsIwEE7is_openEv _ZNKSt13basic_filebufIwSt11char_traitsIwEE7is_openEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv _ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE26_M_destroy_internal_bufferEv _ZNSt13basic_filebufIwSt11char_traitsIwEE26_M_destroy_internal_bufferEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE22_M_convert_to_externalEPwx _ZNSt13basic_filebufIwSt11char_traitsIwEE22_M_convert_to_externalEPwx .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE14_M_get_ext_posERi _ZNSt13basic_filebufIwSt11char_traitsIwEE14_M_get_ext_posERi .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE19_M_terminate_outputEv _ZNSt13basic_filebufIwSt11char_traitsIwEE19_M_terminate_outputEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE7_M_seekExSt12_Ios_Seekdiri _ZNSt13basic_filebufIwSt11char_traitsIwEE7_M_seekExSt12_Ios_Seekdiri .text$_ZNs      St13basic_filebufIwSt11char_traitsIwEE8overflowEt _ZNSt13basic_filebufIwSt11char_traitsIwEE8overflowEt .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt13basic_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode _ZNSt13basic_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE5imbueERKSt6locale _ZNSt13basic_filebufIwSt11char_traitsIwEE5imbueERKSt6locale .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE13_M_set_bufferEx _ZNSt13basic_filebufIwSt11char_traitsIwEE13_M_set_bufferEx .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EOS2_ _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EOS2_ .rdata$_ZTCSt14basic_ifstreamIwSt11char_traitsIwEE0_St13basic_istreamIwS1_E .rdata$_ZTVSt14basic_ifstreamIwSt11cht      ar_traitsIwEE .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt14basic_ifstreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE5rdbufEv _ZNKSt14basic_ifstreamIwSt11char_traitsIwEE5rdbufEv .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv _ZNSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .text$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv _ZNKSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EOS2_ _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EOS2_ .rdata$_ZTCSt14basic_ofstreamIwSt11char_traitsIwEE0_St13basic_ostreamIwS1_E .rdata$_ZTVSt14basic_ofstreamIwSt11char_traitsIwEE .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt14basic_ofstreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNKSt14basic_ofstreamIwSt11char_traitsIwEE5rdbufEv _ZNKSt14basic_ofstreamIwSt11char_traitsIwEE5ru      dbufEv .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv _ZNSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .text$_ZNKSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv _ZNKSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EOS2_ _ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EOS2_ .rdata$_ZTCSt13basic_fstreamIwSt11char_traitsIwEE0_St13basic_istreamIwS1_E .rdata$_ZTVSt13basic_fstreamIwSt11char_traitsIwEE .rdata$_ZTCSt13basic_fstreamIwSt11char_traitsIwEE16_St13basic_ostreamIwS1_E .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt13basic_fstreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNKSt13basic_fstreamIwSt11char_traitsIwEE5rdbufEv _ZNKSt13basic_fstreamIwSt11char_traitsIwEE5rdbufEv .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv _ZNSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .text$_ZNKSt13basic_fstreamIwSt11char_traitsIwv      EE7is_openEv _ZNKSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .text$_ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD1Ev _ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD1Ev .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE5closeEv _ZNSt13basic_filebufIcSt11char_traitsIcEE5closeEv .text$_ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev _ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev .text$_ZNSt13basic_filebufIcSt11char_traitsIcEED1Ev _ZNSt13basic_filebufIcSt11char_traitsIcEED1Ev .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ew      v .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev .text$_ZNSt13basic_filebufIcSt11char_traitsIcEEaSEOS2_ _ZNSt13basic_filebufIcSt11char_traitsIcEEaSEOS2_ .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEaSEOS2_ _ZNSt14basic_ifstreamIcSt11char_traitsIcEEaSEOS2_ .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEaSEOS2_ _ZNSt13basic_fstreamIcSt11char_traitsIcEEaSEOS2_ .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEaSEOS2_ _ZNSt14basic_ofstreamIcSt11char_traitsIcEEaSEOS2_ .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11chx      ar_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNSt13bay      sic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Opez      nmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIcSt1{      1char_traitsIcEE5closeEv _ZNSt14basic_ifstreamIcSt11char_traitsIcEE5closeEv .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv _ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev .text$_ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev _ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev .text$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED1Ev _ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .text$_ZTv0_n2|      4_NSt14basic_ifstreamIcSt11char_traitsIcEED1Ev _ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .text$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .text$_ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev .text$_ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev .text$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .text$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .text$_ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED0Ev _ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .text$_ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev .text$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED0Ev _ZTv0_n}      24_NSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .text$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev .text$_ZZNSt13basic_filebufIwSt11char_traitsIwEE5closeEvEN14__close_sentryD1Ev _ZZNSt13basic_filebufIwSt11char_traitsIwEE5closeEvEN14__close_sentryD1Ev .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE5closeEv _ZNSt13basic_filebufIwSt11char_traitsIwEE5closeEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEED2Ev _ZNSt13basic_filebufIwSt11char_traitsIwEED2Ev .text$_ZNSt13basic_filebufIwSt11char_traitsIwEED1Ev _ZNSt13basic_filebufIwSt11char_traitsIwEED1Ev .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2Ev _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1Ev _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1Ev .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2Ev _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1Ev _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1Ev ~      .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2Ev _ZNSt13basic_fstreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1Ev _ZNSt13basic_fstreamIwSt11char_traitsIwEEC1Ev .text$_ZNSt13basic_filebufIwSt11char_traitsIwEEaSEOS2_ _ZNSt13basic_filebufIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt14basic_ifstreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt13basic_fstreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt14basic_ofstreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode _ZNSt13basic_filebufIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt13basic_filebufIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_      traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11ch�      ar_traitsIwEE4openEPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt13basic_fstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode �      .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode _ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEE�      ESt13_Ios_Openmode _ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE5closeEv _ZNSt14basic_ifstreamIwSt11char_traitsIwEE5closeEv .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE5closeEv _ZNSt14basic_ofstreamIwSt11char_traitsIwEE5closeEv .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEE5closeEv _ZNSt13basic_fstreamIwSt11char_traitsIwEE5closeEv .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED2Ev _ZNSt14basic_ofstreamIwSt11char_traitsIwEED2Ev .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED2Ev _ZNSt14basic_ifstreamIwSt11char_traitsIwEED2Ev .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED1Ev _ZNSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED1Ev _ZNSt14basic_ifstreamIwSt11char_traitsIwEED1Ev .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEED1Ev _ZNSt13basic_fstreamIwSt11char_traitsIwEED1Ev .text$_ZNSt13basic_filebufIwSt11char_traitsIwEED0Ev _ZNSt13basic_filebuf�      IwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .text$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev _ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED1Ev .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEED2Ev _ZNSt13basic_fstreamIwSt11char_traitsIwEED2Ev .text$_ZNSt13basic_fstreamIwSt11char_traitsIwEED0Ev _ZNSt13basic_fstreamIwSt11char_traitsIwEED0Ev .text$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED0Ev _ZNSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .text$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED0Ev _ZNSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSt13b�      asic_fstreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .text$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev _ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .rdata$_ZTSN10__cxxabiv115__forced_unwindE .rdata$_ZTIN10__cxxabiv115__forced_unwindE .rdata$_ZTSSt13basic_filebufIcSt11char_traitsIcEE .rdata$_ZTISt13basic_filebufIcSt11char_traitsIcEE .rdata$_ZTSSt14basic_ifstreamIcSt11char_traitsIcEE .rdata$_ZTISt14basic_ifstreamIcSt11char_traitsIcEE .rdata$_ZTSSt14basic_ofstreamIcSt11char_traitsIcEE .rdata$_ZTISt14basic_ofstreamIcSt11char_traitsIcEE .rdata$_ZTSSt13basic_fstreamIcSt11char_traitsIcEE .rdata$_ZTISt13basic_fstreamIcSt11char_traitsIcEE .rdata$_ZTSSt13basic_filebufIwSt11char_traitsIwEE .rdata$_ZTISt13basic_filebufIwSt11char_traitsIwEE .rdata$_ZTSSt14basic_ifstreamIwSt11char_traitsIwEE .rdata$_ZTISt14basic_ifstreamIwSt11char_traitsIwEE .rdata�      $_ZTSSt14basic_ofstreamIwSt11char_traitsIwEE .rdata$_ZTISt14basic_ofstreamIwSt11char_traitsIwEE .rdata$_ZTSSt13basic_fstreamIwSt11char_traitsIwEE .rdata$_ZTISt13basic_fstreamIwSt11char_traitsIwEE .rdata$_ZTTSt14basic_ifstreamIcSt11char_traitsIcEE .rdata$_ZTTSt14basic_ofstreamIcSt11char_traitsIcEE .rdata$_ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Sd .rdata$_ZTTSt13basic_fstreamIcSt11char_traitsIcEE .rdata$_ZTTSt14basic_ifstreamIwSt11char_traitsIwEE .rdata$_ZTTSt14basic_ofstreamIwSt11char_traitsIwEE .rdata$_ZTCSt13basic_fstreamIwSt11char_traitsIwEE0_St14basic_iostreamIwS1_E .rdata$_ZTTSt13basic_fstreamIwSt11char_traitsIwEE .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcx .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcx .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6setbufEPwx .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6setbufEPwx .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv .xdata$_ZNSt13basic_file�      bufIwSt11char_traitsIwEE9showmanycEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE9showmanycEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4syncEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4syncEv .text$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv.part.41 .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv.part.41 .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv.part.41 .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE9pbackfailEt .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE9pbackfailEt .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE9underflowEv .pda�      ta$_ZNSt13basic_filebufIwSt11char_traitsIwEE9underflowEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcx .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcx .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsputnEPKwx .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsputnEPKwx .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcx .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcx .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsgetnEPwx .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE6xsgetnEPwx .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt13basic_filebufIcSt11char_trai�      tsIcEEC1Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC2EOS2_ .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC2EOS2_ .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC1EOS2_ .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEC1EOS2_ .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv .pdata$_ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcx .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcx .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posERi .pd�      ata$_ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posERi .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE19_M_terminate_outputEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE19_M_terminate_outputEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdiri .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdiri .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcE�      E13_M_set_bufferEx .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE13_M_set_bufferEx .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EOS2_ .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EOS2_ .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EOS2_ .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EOS2_ .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv .pdata$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EOS2_ .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EOS2_ .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EOS2_ .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1E�      OS2_ .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv .pdata$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EOS2_ .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EOS2_ .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EOS2_ .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EOS2_ .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE5rdbufEv .pdata$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE5rdbufEv .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNSt13�      basic_fstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv .pdata$_ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE15_M_create_pbackEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE15_M_create_pbackEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE16_M_destroy_pbackEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE16_M_destroy_pbackEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNKSt13basic_fi�      lebufIwSt11char_traitsIwEE7is_openEv .pdata$_ZNKSt13basic_filebufIwSt11char_traitsIwEE7is_openEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE27_M_allocate_internal_bufferEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE26_M_destroy_internal_bufferEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE26_M_destroy_internal_bufferEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE22_M_convert_to_externalEPwx .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE22_M_convert_to_externalEPwx .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE14_M_get_ext_posERi .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE14_M_get_ext_posERi .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE19_M_terminate_outputEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE19_M_terminate_outputEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7_M_seekExSt12_Ios_Seekdiri .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7_M_seekExSt12_Ios_Seekdiri .xdata$_ZNSt13b�      asic_filebufIwSt11char_traitsIwEE8overflowEt .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE8overflowEt .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE5imbueERKSt6locale .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE5imbueERKSt6locale .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE13_M_set_bufferEx .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE13_M_set_bufferEx .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4swapERS2_ .pd�      ata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE5rdbufEv .pdata$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE5rdbufEv .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNKSt14basic_ifstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNKSt14basic_ofstreamIwSt11char_traitsIwEE5rdbufEv .pdata$_ZNKSt14basic_ofstreamIwSt11char_traitsIwEE5rdbufEv .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZNKSt�      14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNKSt14basic_ofstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNKSt13basic_fstreamIwSt11char_traitsIwEE5rdbufEv .pdata$_ZNKSt13basic_fstreamIwSt11char_traitsIwEE5rdbufEv .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZNKSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .pdata$_ZNKSt13basic_fstreamIwSt11char_traitsIwEE7is_openEv .xdata$_ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD1Ev .pdata$_ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD1Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE5cl�      oseEv .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE5closeEv .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED1Ev .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED1Ev .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ev .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEEaSEOS2_ .pdata$_ZNSt13basic_filebufIcSt11char_tra�      itsIcEEaSEOS2_ .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEaSEOS2_ .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEaSEOS2_ .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEaSEOS2_ .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEaSEOS2_ .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEaSEOS2_ .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEaSEOS2_ .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKNSt7__cx�      x1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char�      _traitsIcEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_�      traitsIcEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKNSt7__cxx1112basic_stringIcS1_SaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIcSt11cha�      r_traitsIcEE5closeEv .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEE5closeEv .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev .xdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev .pdata$_ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev .xdata$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .�      pdata$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED1Ev .xdata$_ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .pdata$_ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED1Ev .xdata$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .pdata$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .xdata$_ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .pdata$_ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev .xdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev .pdata$_ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev .xdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .pdata$_ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .xdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .pdata$_ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .xdata$_ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .pdata$_ZTv0_n24_NSt14basic_ifstreamIcSt11char_traitsIcEED0Ev .xdata$_ZThn16_NSt13basic_fstreamIcSt11�      char_traitsIcEED0Ev .pdata$_ZThn16_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev .xdata$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .pdata$_ZTv0_n24_NSt14basic_ofstreamIcSt11char_traitsIcEED0Ev .xdata$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev .pdata$_ZTv0_n24_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev .xdata$_ZZNSt13basic_filebufIwSt11char_traitsIwEE5closeEvEN14__close_sentryD1Ev .pdata$_ZZNSt13basic_filebufIwSt11char_traitsIwEE5closeEvEN14__close_sentryD1Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE5closeEv .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE5closeEv .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED2Ev .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED2Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED1Ev .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED1Ev .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt14basic_ifstreamIwSt11char_trai�      tsIwEEC1Ev .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4o�      penEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode�       .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE4openEPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt13ba�      sic_fstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1EPKcSt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .�      pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC2ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEEC1ERKNSt7__cxx1112basic_stringIcS0_IcESaIcEEESt13_Ios_Openmode .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE5closeEv .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEE5closeEv .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE5closeEv .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEE5closeEv .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE5closeEv .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEE5closeEv .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED2Ev .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED2Ev .xd�      ata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED2Ev .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED2Ev .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED0Ev .pdata$_ZNSt13basic_filebufIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .xdata$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED1Ev .xdata$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .pdata$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED1Ev .xdata$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEE�      D1Ev .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED2Ev .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED2Ev .xdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt13basic_fstreamIwSt11char_traitsIwEED0Ev .xdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .xdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt14basic_ifstreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt14basic_ofstreamIwSt11char_traitsIwEED0Ev .xdata$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .pdata$_ZThn16_NSt13basic_fstreamIwSt11char_traitsIwEED0Ev .data$.LDFCM0 _ZSt21__throw_bad_exceptionv .rdata$.refptr._ZTVSt13bad_exception .rdata$_ZTISt13�      bad_exception _ZSt17__throw_bad_allocv .rdata$.refptr._ZTVSt9bad_alloc .rdata$_ZTISt9bad_alloc _ZSt16__throw_bad_castv .rdata$.refptr._ZTVSt8bad_cast .rdata$_ZTISt8bad_cast _ZSt18__throw_bad_typeidv .rdata$.refptr._ZTVSt10bad_typeid .rdata$_ZTISt10bad_typeid _ZSt19__throw_logic_errorPKc .rdata$_ZTISt11logic_error _ZSt20__throw_domain_errorPKc .rdata$_ZTISt12domain_error _ZSt24__throw_invalid_argumentPKc .rdata$_ZTISt16invalid_argument _ZSt20__throw_length_errorPKc .rdata$_ZTISt12length_error _ZSt20__throw_out_of_rangePKc .rdata$_ZTISt12out_of_range _ZSt24__throw_out_of_range_fmtPKcz _ZSt21__throw_runtime_errorPKc .rdata$_ZTISt13runtime_error _ZSt19__throw_range_errorPKc .rdata$_ZTISt11range_error _ZSt22__throw_overflow_errorPKc .rdata$_ZTISt14overflow_error _ZSt23__throw_underflow_errorPKc .rdata$_ZTISt15underflow_error .rdata$_ZTSSt13bad_exception .rdata$_ZTSSt8bad_cast .rdata$_ZTSSt10bad_typeid .rdata$_ZTSSt9bad_alloc .rdata$_ZTSSt11logic_error .rdata$_ZTSSt12domain_error .rdata$_ZTSSt16invalid_argu�      ment .rdata$_ZTSSt12length_error .rdata$_ZTSSt12out_of_range .rdata$_ZTSSt13runtime_error .rdata$_ZTSSt11range_error .rdata$_ZTSSt14overflow_error .rdata$_ZTSSt15underflow_error .rdata$.refptr._ZNSt15underflow_errorD1Ev .rdata$.refptr._ZNSt14overflow_errorD1Ev .rdata$.refptr._ZNSt11range_errorD1Ev .rdata$.refptr._ZNSt13runtime_errorD1Ev .rdata$.refptr._ZNSt12out_of_rangeD1Ev .rdata$.refptr._ZNSt12length_errorD1Ev .rdata$.refptr._ZNSt16invalid_argumentD1Ev .rdata$.refptr._ZNSt12domain_errorD1Ev .rdata$.refptr._ZNSt11logic_errorD1Ev .rdata$.refptr._ZNSt10bad_typeidD1Ev .rdata$.refptr._ZNSt8bad_castD1Ev .rdata$.refptr._ZNSt9bad_allocD1Ev .rdata$.refptr._ZNSt13bad_exceptionD1Ev .text$_ZSt21__throw_bad_exceptionv .xdata$_ZSt21__throw_bad_exceptionv .pdata$_ZSt21__throw_bad_exceptionv .text$_ZSt17__throw_bad_allocv .xdata$_ZSt17__throw_bad_allocv .pdata$_ZSt17__throw_bad_allocv .text$_ZSt16__throw_bad_castv .xdata$_ZSt16__throw_bad_castv .pdata$_ZSt16__throw_bad_castv .text$_ZSt18__throw_bad_typeidv .xdata$�      _ZSt18__throw_bad_typeidv .pdata$_ZSt18__throw_bad_typeidv .text$_ZSt19__throw_logic_errorPKc .xdata$_ZSt19__throw_logic_errorPKc .pdata$_ZSt19__throw_logic_errorPKc .text$_ZSt20__throw_domain_errorPKc .xdata$_ZSt20__throw_domain_errorPKc .pdata$_ZSt20__throw_domain_errorPKc .text$_ZSt24__throw_invalid_argumentPKc .xdata$_ZSt24__throw_invalid_argumentPKc .pdata$_ZSt24__throw_invalid_argumentPKc .text$_ZSt20__throw_length_errorPKc .xdata$_ZSt20__throw_length_errorPKc .pdata$_ZSt20__throw_length_errorPKc .text$_ZSt20__throw_out_of_rangePKc .xdata$_ZSt20__throw_out_of_rangePKc .pdata$_ZSt20__throw_out_of_rangePKc .text$_ZSt24__throw_out_of_range_fmtPKcz .xdata$_ZSt24__throw_out_of_range_fmtPKcz .pdata$_ZSt24__throw_out_of_range_fmtPKcz .text$_ZSt21__throw_runtime_errorPKc .xdata$_ZSt21__throw_runtime_errorPKc .pdata$_ZSt21__throw_runtime_errorPKc .text$_ZSt19__throw_range_errorPKc .xdata$_ZSt19__throw_range_errorPKc .pdata$_ZSt19__throw_range_errorPKc .text$_ZSt22__throw_overflow_errorPKc .xdata$_ZSt22__�      throw_overflow_errorPKc .pdata$_ZSt22__throw_overflow_errorPKc .text$_ZSt23__throw_underflow_errorPKc .xdata$_ZSt23__throw_underflow_errorPKc .pdata$_ZSt23__throw_underflow_errorPKc .text$_ZNSt9basic_iosIcSt11char_traitsIcEED1Ev _ZNSt9basic_iosIcSt11char_traitsIcEED1Ev .rdata$_ZTVSt9basic_iosIcSt11char_traitsIcEE .text$_ZNSt9basic_iosIwSt11char_traitsIwEED1Ev _ZNSt9basic_iosIwSt11char_traitsIwEED1Ev .rdata$_ZTVSt9basic_iosIwSt11char_traitsIwEE .text$_ZNSt9basic_iosIcSt11char_traitsIcEED0Ev _ZNSt9basic_iosIcSt11char_traitsIcEED0Ev .text$_ZNSt9basic_iosIwSt11char_traitsIwEED0Ev _ZNSt9basic_iosIwSt11char_traitsIwEED0Ev .text$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvbEv _ZNKSt9basic_iosIcSt11char_traitsIcEEcvbEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEEntEv _ZNKSt9basic_iosIcSt11char_traitsIcEEntEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv _ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv .text$_ZNSt9basic_iosIcSt11char_traitsIcEE5clearESt12_Ios_Iostate _ZNSt9basic_iosIcSt11char_traitsIcEE5clear�      ESt12_Ios_Iostate .text$_ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate _ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate .text$_ZNSt9basic_iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate _ZNSt9basic_iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv _ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv _ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv _ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv _ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv _ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv .text$_ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate _ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate .text$_ZNSt9basic_iosIcSt11char_traitsIcEED2Ev _ZNSt9basic_iosIcSt11char_traitsIcEED2Ev .text$_ZNK�      St9basic_iosIcSt11char_traitsIcEE3tieEv _ZNKSt9basic_iosIcSt11char_traitsIcEE3tieEv .text$_ZNSt9basic_iosIcSt11char_traitsIcEE3tieEPSo _ZNSt9basic_iosIcSt11char_traitsIcEE3tieEPSo .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv _ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv .text$_ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E _ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv _ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv .text$_ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc _ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc _ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc .text$_ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc _ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc .text$_ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev _ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev .text$_ZNSt9basic_iosIcSt11char_traitsIcEEC1Ev _ZNSt9basic_iosIcSt11char_traitsIcEEC1Ev .text$_ZNSt9basic_iosIcSt1�      1char_traitsIcEE9set_rdbufEPSt15basic_streambufIcS1_E _ZNSt9basic_iosIcSt11char_traitsIcEE9set_rdbufEPSt15basic_streambufIcS1_E .text$_ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale _ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale .text$_ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ _ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ .text$_ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale .text$_ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E _ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E .text$_ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E _ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E .text$_ZNSt9basic_iosIcSt11char_traitsIcEEC1EPSt15basic_streambufIcS1_E _ZNSt9basic_iosIcSt11char_traitsIcEEC1EPSt15basic_streambufIcS1_E .text$_ZNSt9basic_iosIcSt11char_traitsIcEE4moveERS2_ _ZNSt9basic_iosIcSt11char_traitsIcEE4moveERS2_ .text$�      _ZNSt9basic_iosIcSt11char_traitsIcEE4swapERS2_ _ZNSt9basic_iosIcSt11char_traitsIcEE4swapERS2_ .text$_ZNSt9basic_iosIcSt11char_traitsIcEE4moveEOS2_ _ZNSt9basic_iosIcSt11char_traitsIcEE4moveEOS2_ .text$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvbEv _ZNKSt9basic_iosIwSt11char_traitsIwEEcvbEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEEntEv _ZNKSt9basic_iosIwSt11char_traitsIwEEntEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE7rdstateEv _ZNKSt9basic_iosIwSt11char_traitsIwEE7rdstateEv .text$_ZNSt9basic_iosIwSt11char_traitsIwEE5clearESt12_Ios_Iostate _ZNSt9basic_iosIwSt11char_traitsIwEE5clearESt12_Ios_Iostate .text$_ZNSt9basic_iosIwSt11char_traitsIwEE8setstateESt12_Ios_Iostate _ZNSt9basic_iosIwSt11char_traitsIwEE8setstateESt12_Ios_Iostate .text$_ZNSt9basic_iosIwSt11char_traitsIwEE11_M_setstateESt12_Ios_Iostate _ZNSt9basic_iosIwSt11char_traitsIwEE11_M_setstateESt12_Ios_Iostate .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE4goodEv _ZNKSt9basic_iosIwSt11char_traitsIwEE4goodEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE3�      eofEv _ZNKSt9basic_iosIwSt11char_traitsIwEE3eofEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE4failEv _ZNKSt9basic_iosIwSt11char_traitsIwEE4failEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE3badEv _ZNKSt9basic_iosIwSt11char_traitsIwEE3badEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE10exceptionsEv _ZNKSt9basic_iosIwSt11char_traitsIwEE10exceptionsEv .text$_ZNSt9basic_iosIwSt11char_traitsIwEE10exceptionsESt12_Ios_Iostate _ZNSt9basic_iosIwSt11char_traitsIwEE10exceptionsESt12_Ios_Iostate .text$_ZNSt9basic_iosIwSt11char_traitsIwEED2Ev _ZNSt9basic_iosIwSt11char_traitsIwEED2Ev .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE3tieEv _ZNKSt9basic_iosIwSt11char_traitsIwEE3tieEv .text$_ZNSt9basic_iosIwSt11char_traitsIwEE3tieEPSt13basic_ostreamIwS1_E _ZNSt9basic_iosIwSt11char_traitsIwEE3tieEPSt13basic_ostreamIwS1_E .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE5rdbufEv _ZNKSt9basic_iosIwSt11char_traitsIwEE5rdbufEv .text$_ZNSt9basic_iosIwSt11char_traitsIwEE5rdbufEPSt15basic_streambufIwS1_E _ZNSt9basic_iosIwSt11char_traitsIw�      EE5rdbufEPSt15basic_streambufIwS1_E .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE4fillEv _ZNKSt9basic_iosIwSt11char_traitsIwEE4fillEv .text$_ZNSt9basic_iosIwSt11char_traitsIwEE4fillEw _ZNSt9basic_iosIwSt11char_traitsIwEE4fillEw .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE6narrowEwc _ZNKSt9basic_iosIwSt11char_traitsIwEE6narrowEwc .text$_ZNKSt9basic_iosIwSt11char_traitsIwEE5widenEc _ZNKSt9basic_iosIwSt11char_traitsIwEE5widenEc .text$_ZNSt9basic_iosIwSt11char_traitsIwEEC2Ev _ZNSt9basic_iosIwSt11char_traitsIwEEC2Ev .text$_ZNSt9basic_iosIwSt11char_traitsIwEEC1Ev _ZNSt9basic_iosIwSt11char_traitsIwEEC1Ev .text$_ZNSt9basic_iosIwSt11char_traitsIwEE9set_rdbufEPSt15basic_streambufIwS1_E _ZNSt9basic_iosIwSt11char_traitsIwEE9set_rdbufEPSt15basic_streambufIwS1_E .text$_ZNSt9basic_iosIwSt11char_traitsIwEE15_M_cache_localeERKSt6locale _ZNSt9basic_iosIwSt11char_traitsIwEE15_M_cache_localeERKSt6locale .text$_ZNSt9basic_iosIwSt11char_traitsIwEE7copyfmtERKS2_ _ZNSt9basic_iosIwSt11char_traitsIwEE7copyfmtERKS2_ .text$_ZNSt9ba�      sic_iosIwSt11char_traitsIwEE5imbueERKSt6locale _ZNSt9basic_iosIwSt11char_traitsIwEE5imbueERKSt6locale .text$_ZNSt9basic_iosIwSt11char_traitsIwEE4initEPSt15basic_streambufIwS1_E _ZNSt9basic_iosIwSt11char_traitsIwEE4initEPSt15basic_streambufIwS1_E .text$_ZNSt9basic_iosIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E _ZNSt9basic_iosIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .text$_ZNSt9basic_iosIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E _ZNSt9basic_iosIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .text$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveERS2_ _ZNSt9basic_iosIwSt11char_traitsIwEE4moveERS2_ .text$_ZNSt9basic_iosIwSt11char_traitsIwEE4swapERS2_ _ZNSt9basic_iosIwSt11char_traitsIwEE4swapERS2_ .text$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveEOS2_ _ZNSt9basic_iosIwSt11char_traitsIwEE4moveEOS2_ .rdata$_ZTSSt8ios_base .rdata$_ZTISt8ios_base .rdata$_ZTSSt9basic_iosIcSt11char_traitsIcEE .rdata$_ZTISt9basic_iosIcSt11char_traitsIcEE .rdata$_ZTSSt9basic_iosIwSt11char_traitsIwEE .rdata$_ZTISt�      9basic_iosIwSt11char_traitsIwEE .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEED1Ev .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEED1Ev .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEED1Ev .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEED1Ev .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEED0Ev .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEED0Ev .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEED0Ev .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEED0Ev .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvbEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvbEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEntEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEntEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5clearESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5clearESt12_Ios_Iostate .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate .xdata$_ZNSt9basic�      _iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEED2Ev .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEED2Ev .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3tieEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE3tieEv .xdata$_ZNSt�      9basic_iosIcSt11char_traitsIcEE3tieEPSo .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE3tieEPSo .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC1Ev .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE9set_rd�      bufEPSt15basic_streambufIcS1_E .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE9set_rdbufEPSt15basic_streambufIcS1_E .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC1EPSt15basic_streambufIcS1_E .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEEC1EPSt15basic_streambufIcS1_E .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4moveERS2_ .pdata$_ZNSt9basic_i�      osIcSt11char_traitsIcEE4moveERS2_ .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4moveEOS2_ .pdata$_ZNSt9basic_iosIcSt11char_traitsIcEE4moveEOS2_ .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvbEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvbEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEntEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEntEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE7rdstateEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE7rdstateEv .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5clearESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5clearESt12_Ios_Iostate .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE8setstateESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE8setstateESt12_Ios_Iostate .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE11_M_setstateESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE11_M_setstateESt12_Ios_Iostate .xdata$_ZNKSt9basic_iosIwSt11char_tr�      aitsIwEE4goodEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE4goodEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3eofEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3eofEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE4failEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE4failEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3badEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3badEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE10exceptionsEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE10exceptionsEv .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE10exceptionsESt12_Ios_Iostate .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE10exceptionsESt12_Ios_Iostate .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEED2Ev .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEED2Ev .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3tieEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE3tieEv .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE3tieEPSt13basic_ostreamIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE3tieEPSt13basic_ostreamIwS1_E .xdata$_ZNKSt9basic_iosIwSt11cha�      r_traitsIwEE5rdbufEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE5rdbufEv .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5rdbufEPSt15basic_streambufIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5rdbufEPSt15basic_streambufIwS1_E .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE4fillEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE4fillEv .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4fillEw .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4fillEw .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE6narrowEwc .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE6narrowEwc .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE5widenEc .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEE5widenEc .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE9set_rdbufEPSt15basic_streambufIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE9set_rdbufEPSt15basic_streambufIwS1_E .xdata$_ZNSt�      9basic_iosIwSt11char_traitsIwEE15_M_cache_localeERKSt6locale .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE15_M_cache_localeERKSt6locale .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE7copyfmtERKS2_ .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE7copyfmtERKS2_ .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5imbueERKSt6locale .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE5imbueERKSt6locale .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4initEPSt15basic_streambufIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4initEPSt15basic_streambufIwS1_E .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveERS2_ .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveERS2_ .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt9basic_iosIwSt11char_tra�      itsIwEE4swapERS2_ .xdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveEOS2_ .pdata$_ZNSt9basic_iosIwSt11char_traitsIwEE4moveEOS2_ _ZNSt8ios_baseC2Ev .rdata$_ZTVSt8ios_base _ZNSt8ios_baseC1Ev _ZNSt8ios_base6xallocEv _ZZNSt8ios_base6xallocEvE6_S_top _ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi _ZNSt8ios_base13_M_grow_wordsEib .rdata$.refptr._ZSt7nothrow _ZNSt8ios_base17_M_call_callbacksENS_5eventE _ZNSt8ios_base20_M_dispose_callbacksEv _ZNSt8ios_baseD2Ev _ZNSt8ios_baseD1Ev _ZNSt8ios_baseD0Ev _ZNSt8ios_base7_M_moveERS_ _ZNSt8ios_base7_M_swapERS_ .text$_ZNSt8ios_baseC2Ev .xdata$_ZNSt8ios_baseC2Ev .pdata$_ZNSt8ios_baseC2Ev .text$_ZNSt8ios_base6xallocEv .xdata$_ZNSt8ios_base6xallocEv .pdata$_ZNSt8ios_base6xallocEv .text$_ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi .xdata$_ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi .pdata$_ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi .text$_ZNSt8ios_base13_M_grow_wordsEib .xdata$_ZNSt8ios_base13_M_grow_wordsEib .pdata$_ZNSt8ios_base13_M_grow_w�      ordsEib .text$_ZNSt8ios_base17_M_call_callbacksENS_5eventE .xdata$_ZNSt8ios_base17_M_call_callbacksENS_5eventE .pdata$_ZNSt8ios_base17_M_call_callbacksENS_5eventE .text$_ZNSt8ios_base20_M_dispose_callbacksEv .xdata$_ZNSt8ios_base20_M_dispose_callbacksEv .pdata$_ZNSt8ios_base20_M_dispose_callbacksEv .text$_ZNSt8ios_baseD2Ev .xdata$_ZNSt8ios_baseD2Ev .pdata$_ZNSt8ios_baseD2Ev .text$_ZNSt8ios_baseD0Ev .xdata$_ZNSt8ios_baseD0Ev .pdata$_ZNSt8ios_baseD0Ev .text$_ZNSt8ios_base7_M_moveERS_ .xdata$_ZNSt8ios_base7_M_moveERS_ .pdata$_ZNSt8ios_base7_M_moveERS_ .text$_ZNSt8ios_base7_M_swapERS_ .xdata$_ZNSt8ios_base7_M_swapERS_ .pdata$_ZNSt8ios_base7_M_swapERS_ .data$_ZZNSt8ios_base6xallocEvE6_S_top .data$_ZNSt8ios_base4Init20_S_synced_with_stdioE .data$_ZNSt8ios_base4Init11_S_refcountE .rdata$_ZNSt8ios_base3endE .rdata$_ZNSt8ios_base3curE .rdata$_ZNSt8ios_base3begE .rdata$_ZNSt8ios_base5truncE .rdata$_ZNSt8ios_base3outE .rdata$_ZNSt8ios_base2inE .rdata$_ZNSt8ios_base6binaryE .rdata$_ZNSt8ios_base3ateE .rdata$_ZNSt�      8ios_base3appE .rdata$_ZNSt8ios_base7goodbitE .rdata$_ZNSt8ios_base7failbitE .rdata$_ZNSt8ios_base6eofbitE .rdata$_ZNSt8ios_base6badbitE .rdata$_ZNSt8ios_base10floatfieldE .rdata$_ZNSt8ios_base9basefieldE .rdata$_ZNSt8ios_base11adjustfieldE .rdata$_ZNSt8ios_base9uppercaseE .rdata$_ZNSt8ios_base7unitbufE .rdata$_ZNSt8ios_base6skipwsE .rdata$_ZNSt8ios_base7showposE .rdata$_ZNSt8ios_base9showpointE .rdata$_ZNSt8ios_base8showbaseE .rdata$_ZNSt8ios_base10scientificE .rdata$_ZNSt8ios_base5rightE .rdata$_ZNSt8ios_base3octE .rdata$_ZNSt8ios_base4leftE .rdata$_ZNSt8ios_base8internalE .rdata$_ZNSt8ios_base3hexE .rdata$_ZNSt8ios_base5fixedE .rdata$_ZNSt8ios_base3decE .rdata$_ZNSt8ios_base9boolalphaE .text$_ZNSdD1Ev _ZNSdD1Ev .rdata$_ZTCSd16_So .rdata$_ZTCSd0_Si .text$_ZNSdD0Ev _ZNSdD0Ev .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEED1Ev _ZNSt14basic_iostreamIwSt11char_traitsIwEED1Ev .rdata$_ZTCSt14basic_iostreamIwSt11char_traitsIwEE16_St13basic_ostreamIwS1_E .rdata$_ZTCSt14basic_iostreamIwSt11char_traitsIwEE0_�      St13basic_istreamIwS1_E .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEED0Ev _ZNSt14basic_iostreamIwSt11char_traitsIwEED0Ev .text$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev _ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSdD1Ev _ZTv0_n24_NSdD1Ev .text$_ZThn16_NSdD1Ev _ZThn16_NSdD1Ev .text$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSdD0Ev _ZTv0_n24_NSdD0Ev .text$_ZThn16_NSdD0Ev _ZThn16_NSdD0Ev .text$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .text$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev _ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .text$_ZSt7setfillIcESt8_SetfillIT_ES1_ _ZSt7setfillIcESt8_SetfillIT_ES1_ .text$_ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSdC1EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSdC1EPSt15basic_streambufIcSt11char_t�      raitsIcEE .rdata$_ZTVSd .text$_ZNSdD2Ev _ZNSdD2Ev .text$_ZNSdC2Ev _ZNSdC2Ev .text$_ZNSdC1Ev _ZNSdC1Ev .text$_ZNSdC2EOSd _ZNSdC2EOSd .text$_ZNSdC1EOSd _ZNSdC1EOSd .text$_ZNSdaSEOSd _ZNSdaSEOSd .text$_ZNSd4swapERSd _ZNSd4swapERSd .text$_ZSt7setfillIwESt8_SetfillIT_ES1_ _ZSt7setfillIwESt8_SetfillIT_ES1_ .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E _ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E _ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .rdata$_ZTVSt14basic_iostreamIwSt11char_traitsIwEE .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEED2Ev _ZNSt14basic_iostreamIwSt11char_traitsIwEED2Ev .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2Ev _ZNSt14basic_iostreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1Ev _ZNSt14basic_iostreamIwSt11char_traitsIwEEC1Ev .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt14�      basic_iostreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EOS2_ _ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EOS2_ .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt14basic_iostreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt14basic_iostreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt14basic_iostreamIwSt11char_traitsIwEE4swapERS2_ .rdata$_ZTSSd .rdata$_ZTISd .rdata$_ZTSSt14basic_iostreamIwSt11char_traitsIwEE .rdata$_ZTISt14basic_iostreamIwSt11char_traitsIwEE .rdata$_ZTTSd .rdata$_ZTTSt14basic_iostreamIwSt11char_traitsIwEE .xdata$_ZNSdD1Ev .pdata$_ZNSdD1Ev .xdata$_ZNSdD0Ev .pdata$_ZNSdD0Ev .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED0Ev .xdata$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .pdata$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .xdata$_ZTv0_n24_NSdD1Ev .pdata$_ZTv0_n24_NSdD1Ev �      .xdata$_ZThn16_NSdD1Ev .pdata$_ZThn16_NSdD1Ev .xdata$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED1Ev .xdata$_ZTv0_n24_NSdD0Ev .pdata$_ZTv0_n24_NSdD0Ev .xdata$_ZThn16_NSdD0Ev .pdata$_ZThn16_NSdD0Ev .xdata$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .xdata$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .pdata$_ZThn16_NSt14basic_iostreamIwSt11char_traitsIwEED0Ev .xdata$_ZSt7setfillIcESt8_SetfillIT_ES1_ .pdata$_ZSt7setfillIcESt8_SetfillIT_ES1_ .xdata$_ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSdC1EPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSdC1EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSdD2Ev .pdata$_ZNSdD2Ev .xdata$_ZNSdC2Ev .pdata$_ZNSdC2Ev .xdata$_ZNSdC1Ev .pdata$_ZNSdC1Ev .xdata$_ZNSdC2EOSd .pdata$_ZNSdC2EOSd .xdata$_ZNSdC1EOSd .pdata$_ZNSdC1EOSd .xdata$_ZNSdaSEOSd�       .pdata$_ZNSdaSEOSd .xdata$_ZNSd4swapERSd .pdata$_ZNSd4swapERSd .xdata$_ZSt7setfillIwESt8_SetfillIT_ES1_ .pdata$_ZSt7setfillIwESt8_SetfillIT_ES1_ .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED2Ev .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEED2Ev .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEC1EOS2_ .x�      data$_ZNSt14basic_iostreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt14basic_iostreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNSiD1Ev _ZNSiD1Ev .rdata$_ZTVSi .text$_ZNSiD0Ev _ZNSiD0Ev .text$_ZNSt13basic_istreamIwSt11char_traitsIwEED1Ev _ZNSt13basic_istreamIwSt11char_traitsIwEED1Ev .rdata$_ZTVSt13basic_istreamIwSt11char_traitsIwEE .text$_ZNSt13basic_istreamIwSt11char_traitsIwEED0Ev _ZNSt13basic_istreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSiD1Ev _ZTv0_n24_NSiD1Ev .text$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSiD0Ev _ZTv0_n24_NSiD0Ev .text$_ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcE�      E _ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSiD2Ev _ZNSiD2Ev .text$_ZNSirsEPFRSiS_E _ZNSirsEPFRSiS_E .text$_ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E _ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .text$_ZNSirsEPFRSt8ios_baseS0_E _ZNSirsEPFRSt8ios_baseS0_E .text$_ZNKSi6gcountEv _ZNKSi6gcountEv .text$_ZNSi7getlineEPcx _ZNSi7getlineEPcx .text$_ZNSiC2Ev _ZNSiC2Ev .text$_ZNSiC1Ev _ZNSiC1Ev .text$_ZNSiC2EOSi _ZNSiC2EOSi .text$_ZNSiC1EOSi _ZNSiC1EOSi .text$_ZNSiaSEOSi _ZNSiaSEOSi .text$_ZNSi4swapERSi _ZNSi4swapERSi .text$_ZNSi6sentryC2ERSib _ZNSi6sentryC2ERSib .text$_ZNSi6sentryC1ERSib _ZNSi6sentryC1ERSib .text$_ZNSirsERs _ZNSirsERs .text$_ZNSirsERi _ZNSirsERi .text$_ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE _ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSi3getEv _ZNSi3getEv .text$_ZNSi3getERc _ZNSi3getERc .text$_ZNSi3getEPcxc _ZNSi3getEPcxc .text$_ZNSi3getEPcx _ZNSi3getEPcx .text$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEEc _ZNSi3getERSt15basic_streambufI�      cSt11char_traitsIcEEc .text$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE _ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSi6ignoreEv _ZNSi6ignoreEv .text$_ZNSi4peekEv _ZNSi4peekEv .text$_ZNSi4readEPcx _ZNSi4readEPcx .text$_ZNSi8readsomeEPcx _ZNSi8readsomeEPcx .text$_ZNSi7putbackEc _ZNSi7putbackEc .text$_ZNSi5ungetEv _ZNSi5ungetEv .text$_ZNSi4syncEv _ZNSi4syncEv .text$_ZNSi5tellgEv _ZNSi5tellgEv .text$_ZNSi5seekgESt4fposIiE _ZNSi5seekgESt4fposIiE .text$_ZNSi5seekgExSt12_Ios_Seekdir _ZNSi5seekgExSt12_Ios_Seekdir .text$_ZNKSi6sentrycvbEv _ZNKSi6sentrycvbEv .text$_ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ _ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_RS3_ _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_RS3_ .text$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh .text$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ra _ZStrsISt11ch�      ar_traitsIcEERSt13basic_istreamIcT_ES5_Ra .text$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph .text$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecision _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecis�      ion .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw .text$_ZNSi10_M_extractItEERSiRT_ _ZNSi10_M_extractItEERSiRT_ .text$_ZNSirsERt _ZNSirsERt .text$_ZNSi10_M_extractIjEERSiRT_ _ZNSi10_M_extractIjEERSiRT_ .text$_ZNSirsERj _ZNSirsERj .text$_ZNSi10_M_extractIlEERSiRT_ _ZNSi10_M_extractIlEERSiRT_ .text$_ZNSirsERl _ZNSirsERl .text$_ZNSi10_M_extractImEERSiRT_ _ZNSi10_M_extractImEERSiRT_ .text$_ZNSirsERm _ZNSirsERm .text$_ZNSi10_M_extractIbEERSiRT_ _ZNSi10_M_extractIbEERSiRT_ .text$_ZNSirsERb _ZNSirsERb .text$_ZNSi10_M_extractIxEERSiRT_ _ZNSi10_M_extractIxEERSiRT_ .text$_ZNSirsERx _ZNSirsERx .text$_ZNSi10_M_extractIyEERSiRT_ _ZNSi10_M_extractIyEERSiRT_ .text$_ZNSirsERy _ZNSirsERy .text$_ZNSi10_M_extractIfEERSiRT_ _ZNSi10_M_extractIfEERSiRT_ .text$_ZNSirsERf _ZNSirsERf .text$_ZNSi10_M_extractIdEERSiRT_ _ZNSi10_M_extractIdEERSiRT_ .text$_ZNSirsERd _ZNSirsERd .text$_ZNSi10_M_extractIeEERSiRT_ _ZNSi10_M_extractIeEERSiRT_ .text$�      _ZNSirsERe _ZNSirsERe .text$_ZNSi10_M_extractIPvEERSiRT_ _ZNSi10_M_extractIPvEERSiRT_ .text$_ZNSirsERPv _ZNSirsERPv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E _ZNSt13basic_istreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E _ZNSt13basic_istreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEED2Ev _ZNSt13basic_istreamIwSt11char_traitsIwEED2Ev .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRS2_S3_E _ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRS2_S3_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt9basic_iosIwS1_ES5_E _ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt9basic_iosIwS1_ES5_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt8ios_baseS4_E _ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt8ios_baseS4_E .text$_ZNKSt13basic_istreamIwSt11char_traitsIwEE6gcountEv _ZNKSt13basic_istreamIwSt11char_traitsIwEE6gcountEv .t�      ext$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwx _ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2Ev _ZNSt13basic_istreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1Ev _ZNSt13basic_istreamIwSt11char_traitsIwEEC1Ev .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt13basic_istreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EOS2_ _ZNSt13basic_istreamIwSt11char_traitsIwEEC1EOS2_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt13basic_istreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt13basic_istreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC2ERS2_b _ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC2ERS2_b .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC1ERS2_b _ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC1ERS2_b .text$_ZNSt13basic_istreamIwSt11char_traitsIwE�      ErsERs _ZNSt13basic_istreamIwSt11char_traitsIwEErsERs .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERi _ZNSt13basic_istreamIwSt11char_traitsIwEErsERi .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPSt15basic_streambufIwS1_E _ZNSt13basic_istreamIwSt11char_traitsIwEErsEPSt15basic_streambufIwS1_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEv _ZNSt13basic_istreamIwSt11char_traitsIwEE3getEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERw _ZNSt13basic_istreamIwSt11char_traitsIwEE3getERw .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwxw _ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwxw .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwx _ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_Ew _ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_Ew .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_E _ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_stre�      ambufIwS1_E .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEv _ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE4peekEv _ZNSt13basic_istreamIwSt11char_traitsIwEE4peekEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE4readEPwx _ZNSt13basic_istreamIwSt11char_traitsIwEE4readEPwx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE8readsomeEPwx _ZNSt13basic_istreamIwSt11char_traitsIwEE8readsomeEPwx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE7putbackEw _ZNSt13basic_istreamIwSt11char_traitsIwEE7putbackEw .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE5ungetEv _ZNSt13basic_istreamIwSt11char_traitsIwEE5ungetEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE4syncEv _ZNSt13basic_istreamIwSt11char_traitsIwEE4syncEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE5tellgEv _ZNSt13basic_istreamIwSt11char_traitsIwEE5tellgEv .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgESt4fposIiE _ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgESt4fposIiE .text$_ZNSt13basic�      _istreamIwSt11char_traitsIwEE5seekgExSt12_Ios_Seekdir _ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgExSt12_Ios_Seekdir .text$_ZNKSt13basic_istreamIwSt11char_traitsIwEE6sentrycvbEv _ZNKSt13basic_istreamIwSt11char_traitsIwEE6sentrycvbEv .text$_ZSt2wsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_ _ZSt2wsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_ .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_RS3_ _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_RS3_ .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_PS3_ _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_PS3_ .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags _ZStrsIwSt11char_traitsIwEER�      St13basic_istreamIT_T0_ES6_St14_Resetiosflags .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_Setbase _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_Setbase .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St13_Setprecision _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St13_Setprecision .text$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St5_Setw _ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St5_Setw .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractItEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractItEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERt _ZNSt13basic_istreamIwSt11char_traitsIwEErsERt .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIjEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIjEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERj _ZNSt13basic_istreamIwSt11char_traitsIwEErsERj .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIlEERS2_RT_ _�      ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIlEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERl _ZNSt13basic_istreamIwSt11char_traitsIwEErsERl .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractImEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractImEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERm _ZNSt13basic_istreamIwSt11char_traitsIwEErsERm .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIbEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIbEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERb _ZNSt13basic_istreamIwSt11char_traitsIwEErsERb .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIxEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIxEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERx _ZNSt13basic_istreamIwSt11char_traitsIwEErsERx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIyEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIyEERS2_RT_ .text$_Z�      NSt13basic_istreamIwSt11char_traitsIwEErsERy _ZNSt13basic_istreamIwSt11char_traitsIwEErsERy .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIfEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIfEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERf _ZNSt13basic_istreamIwSt11char_traitsIwEErsERf .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIdEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIdEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERd _ZNSt13basic_istreamIwSt11char_traitsIwEErsERd .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIeEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIeEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERe _ZNSt13basic_istreamIwSt11char_traitsIwEErsERe .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIPvEERS2_RT_ _ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIPvEERS2_RT_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERPv _ZNSt13basic_istreamIwSt�      11char_traitsIwEErsERPv .rdata$_ZTSSi .rdata$_ZTISi .rdata$_ZTSSt13basic_istreamIwSt11char_traitsIwEE .rdata$_ZTISt13basic_istreamIwSt11char_traitsIwEE .rdata$_ZTTSi .rdata$_ZTTSt13basic_istreamIwSt11char_traitsIwEE .xdata$_ZNSiD1Ev .pdata$_ZNSiD1Ev .xdata$_ZNSiD0Ev .pdata$_ZNSiD0Ev .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSiD1Ev .pdata$_ZTv0_n24_NSiD1Ev .xdata$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED1Ev .xdata$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt13basic_istreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSiD0Ev .pdata$_ZTv0_n24_NSiD0Ev .xdata$_ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcEE .pdat�      a$_ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSiD2Ev .pdata$_ZNSiD2Ev .xdata$_ZNSirsEPFRSiS_E .pdata$_ZNSirsEPFRSiS_E .xdata$_ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .pdata$_ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .xdata$_ZNSirsEPFRSt8ios_baseS0_E .pdata$_ZNSirsEPFRSt8ios_baseS0_E .xdata$_ZNKSi6gcountEv .pdata$_ZNKSi6gcountEv .xdata$_ZNSi7getlineEPcx .pdata$_ZNSi7getlineEPcx .xdata$_ZNSiC2Ev .pdata$_ZNSiC2Ev .xdata$_ZNSiC1Ev .pdata$_ZNSiC1Ev .xdata$_ZNSiC2EOSi .pdata$_ZNSiC2EOSi .xdata$_ZNSiC1EOSi .pdata$_ZNSiC1EOSi .xdata$_ZNSiaSEOSi .pdata$_ZNSiaSEOSi .xdata$_ZNSi4swapERSi .pdata$_ZNSi4swapERSi .xdata$_ZNSi6sentryC2ERSib .pdata$_ZNSi6sentryC2ERSib .xdata$_ZNSi6sentryC1ERSib .pdata$_ZNSi6sentryC1ERSib .xdata$_ZNSirsERs .pdata$_ZNSirsERs .xdata$_ZNSirsERi .pdata$_ZNSirsERi .xdata$_ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSi3getEv .pdata$_ZNSi3getEv .xdata$_ZNSi3getERc .pdata$_ZNSi3getERc .xdata$_�      ZNSi3getEPcxc .pdata$_ZNSi3getEPcxc .xdata$_ZNSi3getEPcx .pdata$_ZNSi3getEPcx .xdata$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEEc .pdata$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEEc .xdata$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSi6ignoreEv .pdata$_ZNSi6ignoreEv .xdata$_ZNSi4peekEv .pdata$_ZNSi4peekEv .xdata$_ZNSi4readEPcx .pdata$_ZNSi4readEPcx .xdata$_ZNSi8readsomeEPcx .pdata$_ZNSi8readsomeEPcx .xdata$_ZNSi7putbackEc .pdata$_ZNSi7putbackEc .xdata$_ZNSi5ungetEv .pdata$_ZNSi5ungetEv .xdata$_ZNSi4syncEv .pdata$_ZNSi4syncEv .xdata$_ZNSi5tellgEv .pdata$_ZNSi5tellgEv .xdata$_ZNSi5seekgESt4fposIiE .pdata$_ZNSi5seekgESt4fposIiE .xdata$_ZNSi5seekgExSt12_Ios_Seekdir .pdata$_ZNSi5seekgExSt12_Ios_Seekdir .xdata$_ZNKSi6sentrycvbEv .pdata$_ZNKSi6sentrycvbEv .xdata$_ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ .pdata$_ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ .xdata$_ZStrsIcSt11char_traitsIcEERS�      t13basic_istreamIT_T0_ES6_RS3_ .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_RS3_ .xdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh .pdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh .xdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ra .pdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ra .xdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph .pdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph .xdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa .pdata$_ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags .pdata$_ZStrsIcSt11char_t�      raitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecision .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecision .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw .xdata$_ZNSi10_M_extractItEERSiRT_ .pdata$_ZNSi10_M_extractItEERSiRT_ .xdata$_ZNSirsERt .pdata$_ZNSirsERt .xdata$_ZNSi10_M_extractIjEERSiRT_ .pdata$_ZNSi10_M_extractIjEERSiRT_ .xdata$_ZNSirsERj .pdata$_ZNSirsERj .xdata$_ZNSi10_M_extractIlEERSiRT_ .pdata$_ZNSi10_M_extractIlEERSiRT_ .xdata$_ZNSirsERl .pdata$_ZNSirsERl .xdata$_ZNSi10_M_extractImEERSiRT_ .pdata$_ZNSi10_M_extractImEERSiRT_ .xdata$_ZNSirsERm .pdata$_ZNSirsERm .xdata$_ZNSi10_M_extractIbEERSiRT_ .pdata$_ZNSi10_M_extractIbEERSiRT_ .xdata$_ZNSirsER�      b .pdata$_ZNSirsERb .xdata$_ZNSi10_M_extractIxEERSiRT_ .pdata$_ZNSi10_M_extractIxEERSiRT_ .xdata$_ZNSirsERx .pdata$_ZNSirsERx .xdata$_ZNSi10_M_extractIyEERSiRT_ .pdata$_ZNSi10_M_extractIyEERSiRT_ .xdata$_ZNSirsERy .pdata$_ZNSirsERy .xdata$_ZNSi10_M_extractIfEERSiRT_ .pdata$_ZNSi10_M_extractIfEERSiRT_ .xdata$_ZNSirsERf .pdata$_ZNSirsERf .xdata$_ZNSi10_M_extractIdEERSiRT_ .pdata$_ZNSi10_M_extractIdEERSiRT_ .xdata$_ZNSirsERd .pdata$_ZNSirsERd .xdata$_ZNSi10_M_extractIeEERSiRT_ .pdata$_ZNSi10_M_extractIeEERSiRT_ .xdata$_ZNSirsERe .pdata$_ZNSirsERe .xdata$_ZNSi10_M_extractIPvEERSiRT_ .pdata$_ZNSi10_M_extractIPvEERSiRT_ .xdata$_ZNSirsERPv .pdata$_ZNSirsERPv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_istreamIwSt11char_traits�      IwEED2Ev .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEED2Ev .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRS2_S3_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRS2_S3_E .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt9basic_iosIwS1_ES5_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt9basic_iosIwS1_ES5_E .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt8ios_baseS4_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPFRSt8ios_baseS4_E .xdata$_ZNKSt13basic_istreamIwSt11char_traitsIwEE6gcountEv .pdata$_ZNKSt13basic_istreamIwSt11char_traitsIwEE6gcountEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt13basic_istreamI�      wSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC2ERS2_b .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC2ERS2_b .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC1ERS2_b .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6sentryC1ERS2_b .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERs .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERs .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERi .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERi .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsEPSt15basic_streambufIwS1_E .xdata$_ZNSt13basi�      c_istreamIwSt11char_traitsIwEE3getEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERw .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERw .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwxw .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwxw .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getEPwx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_Ew .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_Ew .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE3getERSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4peekEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4peekEv .xdata$_ZNSt13basic_istreamIwSt1�      1char_traitsIwEE4readEPwx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4readEPwx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE8readsomeEPwx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE8readsomeEPwx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7putbackEw .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7putbackEw .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5ungetEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5ungetEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4syncEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE4syncEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5tellgEv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5tellgEv .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgESt4fposIiE .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgESt4fposIiE .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgExSt12_Ios_Seekdir .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE5seekgExSt12_Ios_Seekdir .xdata$_ZNKSt13basic_istreamIwSt11char_traitsIwEE6sentrycvbEv .pdata$_ZN�      KSt13basic_istreamIwSt11char_traitsIwEE6sentrycvbEv .xdata$_ZSt2wsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_ .pdata$_ZSt2wsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_ .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_RS3_ .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_RS3_ .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_PS3_ .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_PS3_ .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_Setbase .pdata$_ZStrsIwS�      t11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St8_Setbase .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St13_Setprecision .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St13_Setprecision .xdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St5_Setw .pdata$_ZStrsIwSt11char_traitsIwEERSt13basic_istreamIT_T0_ES6_St5_Setw .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractItEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractItEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERt .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERt .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIjEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIjEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERj .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERj .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIlEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIlEERS2_RT_ .xdata$_�      ZNSt13basic_istreamIwSt11char_traitsIwEErsERl .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERl .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractImEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractImEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERm .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERm .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIbEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIbEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERb .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERb .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIxEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIxEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIyEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIyEERS2_RT_ .xdata$_ZNSt13ba�      sic_istreamIwSt11char_traitsIwEErsERy .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERy .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIfEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIfEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERf .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERf .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIdEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIdEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERd .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERd .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIeEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIeEERS2_RT_ .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERe .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERe .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIPvEERS2_RT_ .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE10_M_extractIPvEERS2_RT_ .xdata$_ZNSt13basic_is�      treamIwSt11char_traitsIwEErsERPv .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEErsERPv .text$_ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv _ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv .text$_ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv _ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv .text$_ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv _ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv .text$_ZNKSt10moneypunctIcLb0EE13do_pos_formatEv _ZNKSt10moneypunctIcLb0EE13do_pos_formatEv .text$_ZNKSt10moneypunctIcLb0EE13do_neg_formatEv _ZNKSt10moneypunctIcLb0EE13do_neg_formatEv .text$_ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv _ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv .text$_ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv _ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv .text$_ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv _ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv .text$_ZNKSt10moneypunctIcLb1EE13do_pos_formatEv _ZNKSt10moneypunctIcLb1EE13do_pos_formatEv .text$_ZNKSt10moneypunctIcLb1EE13do_neg_formatEv _ZNKSt10moneypunctIcLb1�      EE13do_neg_formatEv .text$_ZNSt17moneypunct_bynameIcLb0EED1Ev _ZNSt17moneypunct_bynameIcLb0EED1Ev .rdata$_ZTVSt17moneypunct_bynameIcLb0EE .text$_ZNSt17moneypunct_bynameIcLb1EED1Ev _ZNSt17moneypunct_bynameIcLb1EED1Ev .rdata$_ZTVSt17moneypunct_bynameIcLb1EE .text$_ZNKSt8numpunctIcE16do_decimal_pointEv _ZNKSt8numpunctIcE16do_decimal_pointEv .text$_ZNKSt8numpunctIcE16do_thousands_sepEv _ZNKSt8numpunctIcE16do_thousands_sepEv .text$_ZNSt15numpunct_bynameIcED1Ev _ZNSt15numpunct_bynameIcED1Ev .rdata$_ZTVSt15numpunct_bynameIcE .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .text$_ZNKSt8messagesIcE7do_openERKSsRKSt6locale _ZNKSt8messagesIcE7do_openERKSsRKSt6locale .text$_ZNKSt8messagesIcE8do_closeEi _ZNKSt8messagesIcE8do_closeEi .text$_ZNKSt7collateIcE7do_hashEPKcS2_ _ZNKSt7collateIcE7do_hashEPKcS2_ .text$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt9money_getIcSt19is�      treambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt17__timepunct_cacheIcED1Ev _ZNSt17__timepunct_cacheIcED1Ev .rdata$_ZTVSt17__timepunct_cacheIcE .text$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt8time_putIcSt19ostreamb�      uf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .rdata$_ZTVSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .text$_ZNSt17moneypunct_bynameIcLb0EED0Ev _ZNSt17moneypunct_bynameIcLb0EED0Ev .text$_ZNSt17moneypunct_bynameIcLb1EED0Ev _ZNSt17moneypunct_bynameIcLb1EED0Ev .text$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt15numpunct_bynameIc�      ED0Ev _ZNSt15numpunct_bynameIcED0Ev .text$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt17__timepunct_cacheIcED0Ev _ZNSt17__timepunct_cacheIcED0Ev .text$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .text$_ZNKSt10moneypunctIcLb0EE11do_groupingEv _ZNKSt1�      0moneypunctIcLb0EE11do_groupingEv .text$_ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv _ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv .text$_ZNKSt10moneypunctIcLb0EE16do_positive_signEv _ZNKSt10moneypunctIcLb0EE16do_positive_signEv .text$_ZNKSt10moneypunctIcLb0EE16do_negative_signEv _ZNKSt10moneypunctIcLb0EE16do_negative_signEv .text$_ZNKSt10moneypunctIcLb1EE11do_groupingEv _ZNKSt10moneypunctIcLb1EE11do_groupingEv .text$_ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv _ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv .text$_ZNKSt10moneypunctIcLb1EE16do_positive_signEv _ZNKSt10moneypunctIcLb1EE16do_positive_signEv .text$_ZNKSt10moneypunctIcLb1EE16do_negative_signEv _ZNKSt10moneypunctIcLb1EE16do_negative_signEv .text$_ZNKSt8numpunctIcE11do_groupingEv _ZNKSt8numpunctIcE11do_groupingEv .text$_ZNKSt8numpunctIcE11do_truenameEv _ZNKSt8numpunctIcE11do_truenameEv .text$_ZNKSt8numpunctIcE12do_falsenameEv _ZNKSt8numpunctIcE12do_falsenameEv .text$_ZNSt8messagesIcED1Ev _ZNSt8messagesIcED1Ev .rdata$_ZTVSt8messagesIcE .text$_ZNSt8me�      ssagesIcED0Ev _ZNSt8messagesIcED0Ev .text$_ZNSt7collateIcED1Ev _ZNSt7collateIcED1Ev .rdata$_ZTVSt7collateIcE .text$_ZNSt7collateIcED0Ev _ZNSt7collateIcED0Ev .text$_ZNSt15messages_bynameIcED1Ev _ZNSt15messages_bynameIcED1Ev .text$_ZNSt15messages_bynameIcED0Ev _ZNSt15messages_bynameIcED0Ev .text$_ZNSt14collate_bynameIcED1Ev _ZNSt14collate_bynameIcED1Ev .text$_ZNSt14collate_bynameIcED0Ev _ZNSt14collate_bynameIcED0Ev .text$_ZNSt11__timepunctIcED1Ev _ZNSt11__timepunctIcED1Ev .rdata$_ZTVSt11__timepunctIcE .text$_ZNSt11__timepunctIcED0Ev _ZNSt11__timepunctIcED0Ev .text$_ZNSt14codecvt_bynameIcciED1Ev _ZNSt14codecvt_bynameIcciED1Ev .rdata$_ZTVSt14codecvt_bynameIcciE .text$_ZNSt14codecvt_bynameIcciED0Ev _ZNSt14codecvt_bynameIcciED0Ev _ZNKSt5ctypeIcE5widenEc.part.22 .text$_ZNKSt7collateIcE12do_transformEPKcS2_ _ZNKSt7collateIcE12do_transformEPKcS2_ .text$_ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ _ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ .text$_ZNSt18__moneypunct_cacheIcLb0EEC2Ey _ZNSt18__moneypunct_cacheIcLb0E�      EC2Ey .text$_ZNSt18__moneypunct_cacheIcLb0EEC1Ey _ZNSt18__moneypunct_cacheIcLb0EEC1Ey .text$_ZNSt18__moneypunct_cacheIcLb0EED2Ev _ZNSt18__moneypunct_cacheIcLb0EED2Ev .text$_ZNSt18__moneypunct_cacheIcLb1EEC2Ey _ZNSt18__moneypunct_cacheIcLb1EEC2Ey .text$_ZNSt18__moneypunct_cacheIcLb1EEC1Ey _ZNSt18__moneypunct_cacheIcLb1EEC1Ey .text$_ZNSt18__moneypunct_cacheIcLb1EED2Ev _ZNSt18__moneypunct_cacheIcLb1EED2Ev .text$_ZNSt10moneypunctIcLb0EEC2Ey _ZNSt10moneypunctIcLb0EEC2Ey .rdata$_ZTVSt10moneypunctIcLb0EE .text$_ZNSt10moneypunctIcLb0EEC1Ey _ZNSt10moneypunctIcLb0EEC1Ey .text$_ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy _ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .text$_ZNSt10moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy _ZNSt10moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .text$_ZNSt10moneypunctIcLb0EEC2EPiPKcy _ZNSt10moneypunctIcLb0EEC2EPiPKcy .text$_ZNSt10moneypunctIcLb0EEC1EPiPKcy _ZNSt10moneypunctIcLb0EEC1EPiPKcy .text$_ZNKSt10moneypunctIcLb0EE13decimal_pointEv _ZNK�      St10moneypunctIcLb0EE13decimal_pointEv .text$_ZNKSt10moneypunctIcLb0EE13thousands_sepEv _ZNKSt10moneypunctIcLb0EE13thousands_sepEv .text$_ZNKSt10moneypunctIcLb0EE8groupingEv _ZNKSt10moneypunctIcLb0EE8groupingEv .text$_ZNKSt10moneypunctIcLb0EE11curr_symbolEv _ZNKSt10moneypunctIcLb0EE11curr_symbolEv .text$_ZNKSt10moneypunctIcLb0EE13positive_signEv _ZNKSt10moneypunctIcLb0EE13positive_signEv .text$_ZNKSt10moneypunctIcLb0EE13negative_signEv _ZNKSt10moneypunctIcLb0EE13negative_signEv .text$_ZNKSt10moneypunctIcLb0EE11frac_digitsEv _ZNKSt10moneypunctIcLb0EE11frac_digitsEv .text$_ZNKSt10moneypunctIcLb0EE10pos_formatEv _ZNKSt10moneypunctIcLb0EE10pos_formatEv .text$_ZNKSt10moneypunctIcLb0EE10neg_formatEv _ZNKSt10moneypunctIcLb0EE10neg_formatEv .text$_ZNSt10moneypunctIcLb1EEC2Ey _ZNSt10moneypunctIcLb1EEC2Ey .rdata$_ZTVSt10moneypunctIcLb1EE .text$_ZNSt10moneypunctIcLb1EEC1Ey _ZNSt10moneypunctIcLb1EEC1Ey .text$_ZNSt10moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEy _ZNSt10moneypunctIcLb1EEC2EPSt18__moneypunct_ca�      cheIcLb1EEy .text$_ZNSt10moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy _ZNSt10moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .text$_ZNSt10moneypunctIcLb1EEC2EPiPKcy _ZNSt10moneypunctIcLb1EEC2EPiPKcy .text$_ZNSt10moneypunctIcLb1EEC1EPiPKcy _ZNSt10moneypunctIcLb1EEC1EPiPKcy .text$_ZNKSt10moneypunctIcLb1EE13decimal_pointEv _ZNKSt10moneypunctIcLb1EE13decimal_pointEv .text$_ZNKSt10moneypunctIcLb1EE13thousands_sepEv _ZNKSt10moneypunctIcLb1EE13thousands_sepEv .text$_ZNKSt10moneypunctIcLb1EE8groupingEv _ZNKSt10moneypunctIcLb1EE8groupingEv .text$_ZNKSt10moneypunctIcLb1EE11curr_symbolEv _ZNKSt10moneypunctIcLb1EE11curr_symbolEv .text$_ZNKSt10moneypunctIcLb1EE13positive_signEv _ZNKSt10moneypunctIcLb1EE13positive_signEv .text$_ZNKSt10moneypunctIcLb1EE13negative_signEv _ZNKSt10moneypunctIcLb1EE13negative_signEv .text$_ZNKSt10moneypunctIcLb1EE11frac_digitsEv _ZNKSt10moneypunctIcLb1EE11frac_digitsEv .text$_ZNKSt10moneypunctIcLb1EE10pos_formatEv _ZNKSt10moneypunctIcLb1EE10pos_formatEv .text$_ZNKSt10moneypun�      ctIcLb1EE10neg_formatEv _ZNKSt10moneypunctIcLb1EE10neg_formatEv .text$_ZNSt17moneypunct_bynameIcLb0EEC2EPKcy _ZNSt17moneypunct_bynameIcLb0EEC2EPKcy .text$_ZNSt17moneypunct_bynameIcLb0EEC1EPKcy _ZNSt17moneypunct_bynameIcLb0EEC1EPKcy .text$_ZNSt17moneypunct_bynameIcLb0EEC2ERKSsy _ZNSt17moneypunct_bynameIcLb0EEC2ERKSsy .text$_ZNSt17moneypunct_bynameIcLb0EEC1ERKSsy _ZNSt17moneypunct_bynameIcLb0EEC1ERKSsy .text$_ZNSt17moneypunct_bynameIcLb0EED2Ev _ZNSt17moneypunct_bynameIcLb0EED2Ev .text$_ZNSt17moneypunct_bynameIcLb1EEC2EPKcy _ZNSt17moneypunct_bynameIcLb1EEC2EPKcy .text$_ZNSt17moneypunct_bynameIcLb1EEC1EPKcy _ZNSt17moneypunct_bynameIcLb1EEC1EPKcy .text$_ZNSt17moneypunct_bynameIcLb1EEC2ERKSsy _ZNSt17moneypunct_bynameIcLb1EEC2ERKSsy .text$_ZNSt17moneypunct_bynameIcLb1EEC1ERKSsy _ZNSt17moneypunct_bynameIcLb1EEC1ERKSsy .text$_ZNSt17moneypunct_bynameIcLb1EED2Ev _ZNSt17moneypunct_bynameIcLb1EED2Ev .text$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt9money_getIcSt19istreambuf_iteratorIcS�      t11char_traitsIcEEEC2Ey .text$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traits�      IcEEEC1Ey .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs .text$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt16__numpunct_cacheIcEC2Ey _ZNSt16__numpunct_cacheIcEC2Ey .text$_ZNSt16__numpunct_cacheIcEC1Ey _ZNSt16__numpunct_cacheIcEC1Ey .text$_ZNSt16__numpunct_cacheIcED2Ev _ZNSt16__numpunct_cacheIcED2Ev .text$_ZNSt8numpunctIcEC2Ey _ZNSt8numpunctIcEC2Ey .rdata$_ZTVSt8numpunctIcE .text$_ZNSt8numpunctIcEC1Ey _ZNSt8numpunctIcEC1Ey .text$_ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEy _ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEy .text$_ZNSt8numpunctIcEC1EPSt16__numpunct_cacheIcEy _ZNSt8numpunctIcEC1E�      PSt16__numpunct_cacheIcEy .text$_ZNSt8numpunctIcEC2EPiy _ZNSt8numpunctIcEC2EPiy .text$_ZNSt8numpunctIcEC1EPiy _ZNSt8numpunctIcEC1EPiy .text$_ZNKSt8numpunctIcE13decimal_pointEv _ZNKSt8numpunctIcE13decimal_pointEv .text$_ZNKSt8numpunctIcE13thousands_sepEv _ZNKSt8numpunctIcE13thousands_sepEv .text$_ZNKSt8numpunctIcE8groupingEv _ZNKSt8numpunctIcE8groupingEv .text$_ZNKSt8numpunctIcE8truenameEv _ZNKSt8numpunctIcE8truenameEv .text$_ZNKSt8numpunctIcE9falsenameEv _ZNKSt8numpunctIcE9falsenameEv .text$_ZNSt15numpunct_bynameIcEC2EPKcy _ZNSt15numpunct_bynameIcEC2EPKcy .text$_ZNSt15numpunct_bynameIcEC1EPKcy _ZNSt15numpunct_bynameIcEC1EPKcy .text$_ZNSt15numpunct_bynameIcEC2ERKSsy _ZNSt15numpunct_bynameIcEC2ERKSsy .text$_ZNSt15numpunct_bynameIcEC1ERKSsy _ZNSt15numpunct_bynameIcEC1ERKSsy .text$_ZNSt15numpunct_bynameIcED2Ev _ZNSt15numpunct_bynameIcED2Ev .text$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt7num_getIcSt19istream�      buf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_�      traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .text$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece _ZNKSt7num�      _putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv .text$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt11__timepunctIcEC2Ey _ZNSt11__timepunctIcEC2Ey .text$_ZNSt11__timepunctIcEC1Ey _ZNSt11__timepunctIcEC1Ey .text$_ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEy _ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEy .text$_ZNSt11__timepunctIcEC1EPSt17__timepunct_cacheIcEy _ZNSt11__timepunctIcEC1EPSt17__timepunct_cacheIcEy .text$_ZNSt11__timepunctIcEC2EPiPKcy _ZNSt11__timepunctIcEC2EPiPKcy .text$_ZNSt11__timepunctIcEC1EPiPKcy _ZNSt11__timepunctIcEC1EPiPKcy .text$_ZNKSt11__timepunctIcE15_M_date_formatsEPPKc _ZNKSt11__timepunctIcE15_M_date_formatsEPPKc .text$_ZNKSt11__timepunctIcE15_M_time_formatsEPPKc _ZNKSt11__tim�      epunctIcE15_M_time_formatsEPPKc .text$_ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc _ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc .text$_ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc _ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc .text$_ZNKSt11__timepunctIcE8_M_am_pmEPPKc _ZNKSt11__timepunctIcE8_M_am_pmEPPKc .text$_ZNKSt11__timepunctIcE7_M_daysEPPKc _ZNKSt11__timepunctIcE7_M_daysEPPKc .text$_ZNKSt11__timepunctIcE19_M_days_abbreviatedEPPKc _ZNKSt11__timepunctIcE19_M_days_abbreviatedEPPKc .text$_ZNKSt11__timepunctIcE9_M_monthsEPPKc _ZNKSt11__timepunctIcE9_M_monthsEPPKc .text$_ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc _ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc .text$_ZNSt11__timepunctIcED2Ev _ZNSt11__timepunctIcED2Ev .text$_ZNSt17__timepunct_cacheIcEC2Ey _ZNSt17__timepunct_cacheIcEC2Ey .text$_ZNSt17__timepunct_cacheIcEC1Ey _ZNSt17__timepunct_cacheIcEC1Ey .text$_ZNSt17__timepunct_cacheIcED2Ev _ZNSt17__timepunct_cacheIcED2Ev .text$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIc�      EEEC2Ey _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc .text$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .rdata$_ZTVSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERK�      Ssy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .text$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .text$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8g�      et_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt8time_getIcSt19is�      treambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .rdata$_ZTVSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .text$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .text$_ZNSt8messagesIcEC2Ey _Z�      NSt8messagesIcEC2Ey .text$_ZNSt8messagesIcEC1Ey _ZNSt8messagesIcEC1Ey .text$_ZNSt8messagesIcEC2EPiPKcy _ZNSt8messagesIcEC2EPiPKcy .text$_ZNSt8messagesIcEC1EPiPKcy _ZNSt8messagesIcEC1EPiPKcy .text$_ZNKSt8messagesIcE4openERKSsRKSt6locale _ZNKSt8messagesIcE4openERKSsRKSt6locale .text$_ZNKSt8messagesIcE4openERKSsRKSt6localePKc _ZNKSt8messagesIcE4openERKSsRKSt6localePKc .text$_ZNKSt8messagesIcE3getEiiiRKSs _ZNKSt8messagesIcE3getEiiiRKSs .text$_ZNKSt8messagesIcE5closeEi _ZNKSt8messagesIcE5closeEi .text$_ZNSt8messagesIcED2Ev _ZNSt8messagesIcED2Ev .text$_ZNKSt8messagesIcE18_M_convert_to_charERKSs _ZNKSt8messagesIcE18_M_convert_to_charERKSs .text$_ZNKSt8messagesIcE20_M_convert_from_charEPc _ZNKSt8messagesIcE20_M_convert_from_charEPc .text$_ZNSt15messages_bynameIcEC2EPKcy _ZNSt15messages_bynameIcEC2EPKcy .rdata$_ZTVSt15messages_bynameIcE .text$_ZNSt15messages_bynameIcEC1EPKcy _ZNSt15messages_bynameIcEC1EPKcy .text$_ZNSt15messages_bynameIcEC2ERKSsy _ZNSt15messages_bynameIcEC2ERKSsy .text$_ZNSt15messages_bynameIc�      EC1ERKSsy _ZNSt15messages_bynameIcEC1ERKSsy .text$_ZNSt15messages_bynameIcED2Ev _ZNSt15messages_bynameIcED2Ev _ZNSt12ctype_bynameIcEC2ERKSsy _ZNSt12ctype_bynameIcEC1ERKSsy .text$_ZNSt14codecvt_bynameIcciEC2EPKcy _ZNSt14codecvt_bynameIcciEC2EPKcy .text$_ZNSt14codecvt_bynameIcciEC1EPKcy _ZNSt14codecvt_bynameIcciEC1EPKcy .text$_ZNSt14codecvt_bynameIcciEC2ERKSsy _ZNSt14codecvt_bynameIcciEC2ERKSsy .text$_ZNSt14codecvt_bynameIcciEC1ERKSsy _ZNSt14codecvt_bynameIcciEC1ERKSsy .text$_ZNSt14codecvt_bynameIcciED2Ev _ZNSt14codecvt_bynameIcciED2Ev .text$_ZNSt7collateIcEC2Ey _ZNSt7collateIcEC2Ey .text$_ZNSt7collateIcEC1Ey _ZNSt7collateIcEC1Ey .text$_ZNSt7collateIcEC2EPiy _ZNSt7collateIcEC2EPiy .text$_ZNSt7collateIcEC1EPiy _ZNSt7collateIcEC1EPiy .text$_ZNKSt7collateIcE7compareEPKcS2_S2_S2_ _ZNKSt7collateIcE7compareEPKcS2_S2_S2_ .text$_ZNKSt7collateIcE9transformEPKcS2_ _ZNKSt7collateIcE9transformEPKcS2_ .text$_ZNKSt7collateIcE4hashEPKcS2_ _ZNKSt7collateIcE4hashEPKcS2_ .text$_ZNSt7collateIcED2Ev _ZNSt7collateIcED2Ev .t�      ext$_ZNSt14collate_bynameIcEC2EPKcy _ZNSt14collate_bynameIcEC2EPKcy .rdata$_ZTVSt14collate_bynameIcE .text$_ZNSt14collate_bynameIcEC1EPKcy _ZNSt14collate_bynameIcEC1EPKcy .text$_ZNSt14collate_bynameIcEC2ERKSsy _ZNSt14collate_bynameIcEC2ERKSsy .text$_ZNSt14collate_bynameIcEC1ERKSsy _ZNSt14collate_bynameIcEC1ERKSsy .text$_ZNSt14collate_bynameIcED2Ev _ZNSt14collate_bynameIcED2Ev .text$_ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale _ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale .text$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt�      12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZSt9use_facetISt7codecvtIcciEERKT_RKSt6locale _ZSt9use_facetISt7codecvtIcciEERKT_RKSt6locale .rdata$_ZTISt7codecvtIcciE .text$_ZSt9use_facetISt7collateIcEERKT_RKSt6locale _ZSt9use_facetISt7collateIcEERKT_RKSt6locale .data$_ZNSt7collateIcE2idE .rdata$_ZTISt7collateIcE .text$_ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale _ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale .data$_ZNSt8numpunctIcE2idE .rdata$_ZTISt8numpunctIcE .text$_ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale _ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt7num_�      getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt10moneypunctIcLb1EEERKT_RKSt6locale _ZSt9use_facetISt10moneypunctIcLb1EEERKT_RKSt6locale .data$_ZNSt10moneypunctIcLb1EE2idE .rdata$_ZTISt10moneypunctIcLb1EE .text$_ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale _ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale _ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale .data$_ZNSt10moneypunctIcLb0EE2idE .rdata$_ZTISt10moneypunctIcLb0EE .text$_ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale _ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt9money_putIcSt19os�      treambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale _ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale .data$_ZNSt11__timepunctIcE2idE .rdata$_ZTISt11__timepunctIcE .text$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc .text$_ZSt9use_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt8time_put�      IcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .data$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .rdata$_ZTISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .text$_ZSt9use_facetISt8messagesIcEERKT_RKSt6locale _ZSt9use_facetISt8messagesIcEERKT_RKSt6locale .data$_ZNSt8messagesIcE2idE .rdata$_ZTISt8messagesIcE .text$_ZSt9has_facetISt5ctypeIcEEbRKSt6locale _ZSt9has_facetISt5ctypeIcEEbRKSt6locale .text$_ZSt9has_facetISt7codecvtIcciEEbRKSt6locale _ZSt9has_facetISt7codecvtIcciEEbRKSt6locale .text$_ZSt9has_facetISt7collateIcEEbRKSt6locale _ZSt9has_facetISt7collateIcEEbRKSt6locale .text$_ZSt9has_facetISt8numpunctIcEEbRKSt6locale _ZSt9has_fa�      cetISt8numpunctIcEEbRKSt6locale .text$_ZSt9has_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale _ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale .text$_ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt11__timepunctIcEEbRKSt6locale _ZSt9has_facetISt11__timepunctIcEEbRKSt6locale .text$_ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorI�      cSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .text$_ZSt9has_facetISt8messagesIcEEbRKSt6locale _ZSt9has_facetISt8messagesIcEEbRKSt6locale .text$_ZSt14__add_groupingIcEPT_S1_S0_PKcyPKS0_S5_ _ZSt14__add_groupingIcEPT_S1_S0_PKcyPKS0_S5_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcycS6_PcS7_Ri _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcycS6_PcS7_Ri .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcycRSt8ios_basePcS9_Ri _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcycRSt8ios_basePcS9_Ri .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs _ZNKSt9money_p�      utIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece .text$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs .text$_ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcxx _ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcxx .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6_M_padEcxRSt8ios_basePcPKcRi _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6_M_padEcxRSt8ios_basePcPKcRi .text$_ZSt13__int_�      to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZSt13__int_to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .text$_ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .text$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale .text$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecl _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_trai�      tsIcEEE3putES3_RSt8ios_basecl .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_RSt8ios_basecT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_RSt8ios_basecT_ .text$_ZNKSt7num_putIcSt19ostrea�      mbuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy _ZNKSt7num_putIcSt19ostreambuf�      _iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ .text$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIcSt19istreambuf_iteratorI�      cSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc _ZNKSt8time_getIcSt19istreambuf_itera�      torIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP�      2tmcc .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_ba�      seRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_�      S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3�      _S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE       14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcS      t11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .text$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNK      St9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSC_ _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSC_ _GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKSsy .data$_ZGVNSt10moneypunctIcLb0EE2idE .data$_ZGVNSt10moneypunctIcLb1EE2idE .data$_ZGVNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt8numpunctIcE2idE .data$_ZGVNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .dat      a$_ZGVNSt11__timepunctIcE2idE .data$_ZGVNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .data$_ZGVNSt8messagesIcE2idE .data$_ZGVNSt7collateIcE2idE .rdata$_ZTSSt7collateIcE .rdata$_ZTSSt14collate_bynameIcE .rdata$_ZTISt14collate_bynameIcE .rdata$_ZTSSt8numpunctIcE .rdata$_ZTSSt15numpunct_bynameIcE .rdata$_ZTISt15numpunct_bynameIcE .rdata$_ZTSSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt17__timepunct_cacheIcE .rdata$_ZTISt17__timepunct_cacheIcE .rdata$_ZTSSt11__timepunctIcE .rdata$_ZTSSt10moneypunctIcLb1EE .rdata$_ZTSSt10moneypunctIcLb0EE .rdata$_ZTSSt8messagesIcE .rdata$_ZTSSt23__codecvt_abstract_baseIcciE .rdata$_ZTISt23__codecvt_abstract_baseIcciE .rdata$_ZTSSt7codecvtIcciE .rdata$_ZTSSt14codecvt_bynameIcciE .rdata$_ZTISt14codecvt_bynameIcciE .rdata$_ZTSSt17moneypunct_bynameIcLb0EE .rdata$_ZTISt17moneypunct_bynameIcLb0      EE .rdata$_ZTSSt17moneypunct_bynameIcLb1EE .rdata$_ZTISt17moneypunct_bynameIcLb1EE .rdata$_ZTSSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTISt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTISt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .rdata$_ZTSSt15messages_bynameIcE .rdata$_ZTISt15messages_bynameIcE .rdata$_ZTSSt21__ctype_abstract_baseIcE .rdata$_ZTISt21__ctype_abstract_baseIcE .rdata$_ZTVSt23__codecvt_abstract_baseIcciE .rdata$_ZTVSt21__ctype_abstract_baseIcE .rdata$_ZNSt17moneypunct_bynameIcLb1EE4intlE .rdata$_ZNSt17moneypunct_bynameIcLb0EE4intlE .rdata$_ZNSt10mon      eypunctIcLb1EE4intlE .rdata$_ZNSt10moneypunctIcLb0EE4intlE .xdata$_ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv .pdata$_ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv .xdata$_ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv .pdata$_ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv .xdata$_ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv .pdata$_ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv .xdata$_ZNKSt10moneypunctIcLb0EE13do_pos_formatEv .pdata$_ZNKSt10moneypunctIcLb0EE13do_pos_formatEv .xdata$_ZNKSt10moneypunctIcLb0EE13do_neg_formatEv .pdata$_ZNKSt10moneypunctIcLb0EE13do_neg_formatEv .xdata$_ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv .pdata$_ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv .xdata$_ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv .pdata$_ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv .xdata$_ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv .pdata$_ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv .xdata$_ZNKSt10moneypunctIcLb1EE13do_pos_formatEv .pdata$_ZNKSt10moneypunctIcLb1EE13do_pos_formatEv .xdata$_ZNKSt10moneypunctIcLb      1EE13do_neg_formatEv .pdata$_ZNKSt10moneypunctIcLb1EE13do_neg_formatEv .xdata$_ZNSt17moneypunct_bynameIcLb0EED1Ev .pdata$_ZNSt17moneypunct_bynameIcLb0EED1Ev .xdata$_ZNSt17moneypunct_bynameIcLb1EED1Ev .pdata$_ZNSt17moneypunct_bynameIcLb1EED1Ev .xdata$_ZNKSt8numpunctIcE16do_decimal_pointEv .pdata$_ZNKSt8numpunctIcE16do_decimal_pointEv .xdata$_ZNKSt8numpunctIcE16do_thousands_sepEv .pdata$_ZNKSt8numpunctIcE16do_thousands_sepEv .xdata$_ZNSt15numpunct_bynameIcED1Ev .pdata$_ZNSt15numpunct_bynameIcED1Ev .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv .xdata$_ZNKSt8messagesIcE7do_openERKSsRKSt6locale .pdata$_ZNKSt8messagesIcE7do_openERKSsRKSt6locale .xdata$_ZNKSt8messagesIcE8do_closeEi .pdata$_ZNKSt8messagesIcE8do_closeEi .xdata$_ZNKSt7collateIcE7do_hashEPKcS2_ .pdata$_ZNKSt7collateIcE7do_hashEPKcS2_ .xdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt9      money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt17__timepunct_cacheIcED1Ev .pdata$_ZNSt17__timepunct_cacheIcED1Ev .xdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_tra      itsIcEEED1Ev .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev .xdata$_ZNSt17moneypunct_bynameIcLb0EED0Ev .pdata$_ZNSt17moneypunct_bynameIcLb0EED0Ev .xdata$_ZNSt17moneypunct_bynameIcLb1EED0Ev .pdata$_ZNSt17moneypunct_bynameIcLb1EED0Ev .xdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt15numpunct_bynameIcED0Ev .pdata$_ZNSt15numpunct_bynameIcED0Ev .xdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNS	      t17__timepunct_cacheIcED0Ev .pdata$_ZNSt17__timepunct_cacheIcED0Ev .xdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev .xdata$_ZNKSt10moneypunctIcLb0EE11do_groupingEv .pdata$_ZNKSt10moneypunctIcLb0EE11do_groupingEv .xdata$_ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv .pdata$_ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv .xdata$_ZNKSt10moneypunctIcLb0EE16do_positive_signEv .pdata$_ZNKSt10moneypunctIcLb0EE16do_positive_signEv .xdata$_ZNKSt10moneypunctIcLb
      0EE16do_negative_signEv .pdata$_ZNKSt10moneypunctIcLb0EE16do_negative_signEv .xdata$_ZNKSt10moneypunctIcLb1EE11do_groupingEv .pdata$_ZNKSt10moneypunctIcLb1EE11do_groupingEv .xdata$_ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv .pdata$_ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv .xdata$_ZNKSt10moneypunctIcLb1EE16do_positive_signEv .pdata$_ZNKSt10moneypunctIcLb1EE16do_positive_signEv .xdata$_ZNKSt10moneypunctIcLb1EE16do_negative_signEv .pdata$_ZNKSt10moneypunctIcLb1EE16do_negative_signEv .xdata$_ZNKSt8numpunctIcE11do_groupingEv .pdata$_ZNKSt8numpunctIcE11do_groupingEv .xdata$_ZNKSt8numpunctIcE11do_truenameEv .pdata$_ZNKSt8numpunctIcE11do_truenameEv .xdata$_ZNKSt8numpunctIcE12do_falsenameEv .pdata$_ZNKSt8numpunctIcE12do_falsenameEv .xdata$_ZNSt8messagesIcED1Ev .pdata$_ZNSt8messagesIcED1Ev .xdata$_ZNSt8messagesIcED0Ev .pdata$_ZNSt8messagesIcED0Ev .xdata$_ZNSt7collateIcED1Ev .pdata$_ZNSt7collateIcED1Ev .xdata$_ZNSt7collateIcED0Ev .pdata$_ZNSt7collateIcED0Ev .xdata$_ZNSt15messages_bynameIcED1Ev .pdata$_ZNSt15me      ssages_bynameIcED1Ev .xdata$_ZNSt15messages_bynameIcED0Ev .pdata$_ZNSt15messages_bynameIcED0Ev .xdata$_ZNSt14collate_bynameIcED1Ev .pdata$_ZNSt14collate_bynameIcED1Ev .xdata$_ZNSt14collate_bynameIcED0Ev .pdata$_ZNSt14collate_bynameIcED0Ev .xdata$_ZNSt11__timepunctIcED1Ev .pdata$_ZNSt11__timepunctIcED1Ev .xdata$_ZNSt11__timepunctIcED0Ev .pdata$_ZNSt11__timepunctIcED0Ev .xdata$_ZNSt14codecvt_bynameIcciED1Ev .pdata$_ZNSt14codecvt_bynameIcciED1Ev .xdata$_ZNSt14codecvt_bynameIcciED0Ev .pdata$_ZNSt14codecvt_bynameIcciED0Ev .text$_ZNKSt5ctypeIcE5widenEc.part.22 .xdata$_ZNKSt5ctypeIcE5widenEc.part.22 .pdata$_ZNKSt5ctypeIcE5widenEc.part.22 .xdata$_ZNKSt7collateIcE12do_transformEPKcS2_ .pdata$_ZNKSt7collateIcE12do_transformEPKcS2_ .xdata$_ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ .pdata$_ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ .xdata$_ZNSt18__moneypunct_cacheIcLb0EEC2Ey .pdata$_ZNSt18__moneypunct_cacheIcLb0EEC2Ey .xdata$_ZNSt18__moneypunct_cacheIcLb0EEC1Ey .pdata$_ZNSt18__moneypunct_cacheIcLb0EEC1Ey .xdata$_Z      NSt18__moneypunct_cacheIcLb0EED2Ev .pdata$_ZNSt18__moneypunct_cacheIcLb0EED2Ev .xdata$_ZNSt18__moneypunct_cacheIcLb1EEC2Ey .pdata$_ZNSt18__moneypunct_cacheIcLb1EEC2Ey .xdata$_ZNSt18__moneypunct_cacheIcLb1EEC1Ey .pdata$_ZNSt18__moneypunct_cacheIcLb1EEC1Ey .xdata$_ZNSt18__moneypunct_cacheIcLb1EED2Ev .pdata$_ZNSt18__moneypunct_cacheIcLb1EED2Ev .xdata$_ZNSt10moneypunctIcLb0EEC2Ey .pdata$_ZNSt10moneypunctIcLb0EEC2Ey .xdata$_ZNSt10moneypunctIcLb0EEC1Ey .pdata$_ZNSt10moneypunctIcLb0EEC1Ey .xdata$_ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .pdata$_ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEy .xdata$_ZNSt10moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .pdata$_ZNSt10moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEy .xdata$_ZNSt10moneypunctIcLb0EEC2EPiPKcy .pdata$_ZNSt10moneypunctIcLb0EEC2EPiPKcy .xdata$_ZNSt10moneypunctIcLb0EEC1EPiPKcy .pdata$_ZNSt10moneypunctIcLb0EEC1EPiPKcy .xdata$_ZNKSt10moneypunctIcLb0EE13decimal_pointEv .pdata$_ZNKSt10moneypunctIcLb0EE13decimal_pointEv .      xdata$_ZNKSt10moneypunctIcLb0EE13thousands_sepEv .pdata$_ZNKSt10moneypunctIcLb0EE13thousands_sepEv .xdata$_ZNKSt10moneypunctIcLb0EE8groupingEv .pdata$_ZNKSt10moneypunctIcLb0EE8groupingEv .xdata$_ZNKSt10moneypunctIcLb0EE11curr_symbolEv .pdata$_ZNKSt10moneypunctIcLb0EE11curr_symbolEv .xdata$_ZNKSt10moneypunctIcLb0EE13positive_signEv .pdata$_ZNKSt10moneypunctIcLb0EE13positive_signEv .xdata$_ZNKSt10moneypunctIcLb0EE13negative_signEv .pdata$_ZNKSt10moneypunctIcLb0EE13negative_signEv .xdata$_ZNKSt10moneypunctIcLb0EE11frac_digitsEv .pdata$_ZNKSt10moneypunctIcLb0EE11frac_digitsEv .xdata$_ZNKSt10moneypunctIcLb0EE10pos_formatEv .pdata$_ZNKSt10moneypunctIcLb0EE10pos_formatEv .xdata$_ZNKSt10moneypunctIcLb0EE10neg_formatEv .pdata$_ZNKSt10moneypunctIcLb0EE10neg_formatEv .xdata$_ZNSt10moneypunctIcLb1EEC2Ey .pdata$_ZNSt10moneypunctIcLb1EEC2Ey .xdata$_ZNSt10moneypunctIcLb1EEC1Ey .pdata$_ZNSt10moneypunctIcLb1EEC1Ey .xdata$_ZNSt10moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEy .pdata$_ZNSt10moneypunctIcLb1EEC2EPSt18      __moneypunct_cacheIcLb1EEy .xdata$_ZNSt10moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .pdata$_ZNSt10moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEy .xdata$_ZNSt10moneypunctIcLb1EEC2EPiPKcy .pdata$_ZNSt10moneypunctIcLb1EEC2EPiPKcy .xdata$_ZNSt10moneypunctIcLb1EEC1EPiPKcy .pdata$_ZNSt10moneypunctIcLb1EEC1EPiPKcy .xdata$_ZNKSt10moneypunctIcLb1EE13decimal_pointEv .pdata$_ZNKSt10moneypunctIcLb1EE13decimal_pointEv .xdata$_ZNKSt10moneypunctIcLb1EE13thousands_sepEv .pdata$_ZNKSt10moneypunctIcLb1EE13thousands_sepEv .xdata$_ZNKSt10moneypunctIcLb1EE8groupingEv .pdata$_ZNKSt10moneypunctIcLb1EE8groupingEv .xdata$_ZNKSt10moneypunctIcLb1EE11curr_symbolEv .pdata$_ZNKSt10moneypunctIcLb1EE11curr_symbolEv .xdata$_ZNKSt10moneypunctIcLb1EE13positive_signEv .pdata$_ZNKSt10moneypunctIcLb1EE13positive_signEv .xdata$_ZNKSt10moneypunctIcLb1EE13negative_signEv .pdata$_ZNKSt10moneypunctIcLb1EE13negative_signEv .xdata$_ZNKSt10moneypunctIcLb1EE11frac_digitsEv .pdata$_ZNKSt10moneypunctIcLb1EE11frac_digitsEv .xdata$_ZNKSt      10moneypunctIcLb1EE10pos_formatEv .pdata$_ZNKSt10moneypunctIcLb1EE10pos_formatEv .xdata$_ZNKSt10moneypunctIcLb1EE10neg_formatEv .pdata$_ZNKSt10moneypunctIcLb1EE10neg_formatEv .xdata$_ZNSt17moneypunct_bynameIcLb0EEC2EPKcy .pdata$_ZNSt17moneypunct_bynameIcLb0EEC2EPKcy .xdata$_ZNSt17moneypunct_bynameIcLb0EEC1EPKcy .pdata$_ZNSt17moneypunct_bynameIcLb0EEC1EPKcy .xdata$_ZNSt17moneypunct_bynameIcLb0EEC2ERKSsy .pdata$_ZNSt17moneypunct_bynameIcLb0EEC2ERKSsy .xdata$_ZNSt17moneypunct_bynameIcLb0EEC1ERKSsy .pdata$_ZNSt17moneypunct_bynameIcLb0EEC1ERKSsy .xdata$_ZNSt17moneypunct_bynameIcLb0EED2Ev .pdata$_ZNSt17moneypunct_bynameIcLb0EED2Ev .xdata$_ZNSt17moneypunct_bynameIcLb1EEC2EPKcy .pdata$_ZNSt17moneypunct_bynameIcLb1EEC2EPKcy .xdata$_ZNSt17moneypunct_bynameIcLb1EEC1EPKcy .pdata$_ZNSt17moneypunct_bynameIcLb1EEC1EPKcy .xdata$_ZNSt17moneypunct_bynameIcLb1EEC2ERKSsy .pdata$_ZNSt17moneypunct_bynameIcLb1EEC2ERKSsy .xdata$_ZNSt17moneypunct_bynameIcLb1EEC1ERKSsy .pdata$_ZNSt17moneypunct_bynameIcLb1EEC1ERKSsy .xdata$_ZNS      t17moneypunct_bynameIcLb1EED2Ev .pdata$_ZNSt17moneypunct_bynameIcLb1EED2Ev .xdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt9money_putIcSt19ostreambuf_      iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece .pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs .pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs .xdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt16__numpunct_cacheIcEC2Ey .pdata$_ZNSt16__numpunct_cacheIcEC2Ey .xdata$_ZNSt16__numpunct_cacheIcEC1Ey .pdata$_ZNSt16__numpunct_cacheIcEC1Ey .xdata$_ZNSt16__numpunct_cacheIcED2Ev .pdata$_ZNSt16__numpunct_cacheIcED2Ev .      xdata$_ZNSt8numpunctIcEC2Ey .pdata$_ZNSt8numpunctIcEC2Ey .xdata$_ZNSt8numpunctIcEC1Ey .pdata$_ZNSt8numpunctIcEC1Ey .xdata$_ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEy .pdata$_ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEy .xdata$_ZNSt8numpunctIcEC1EPSt16__numpunct_cacheIcEy .pdata$_ZNSt8numpunctIcEC1EPSt16__numpunct_cacheIcEy .xdata$_ZNSt8numpunctIcEC2EPiy .pdata$_ZNSt8numpunctIcEC2EPiy .xdata$_ZNSt8numpunctIcEC1EPiy .pdata$_ZNSt8numpunctIcEC1EPiy .xdata$_ZNKSt8numpunctIcE13decimal_pointEv .pdata$_ZNKSt8numpunctIcE13decimal_pointEv .xdata$_ZNKSt8numpunctIcE13thousands_sepEv .pdata$_ZNKSt8numpunctIcE13thousands_sepEv .xdata$_ZNKSt8numpunctIcE8groupingEv .pdata$_ZNKSt8numpunctIcE8groupingEv .xdata$_ZNKSt8numpunctIcE8truenameEv .pdata$_ZNKSt8numpunctIcE8truenameEv .xdata$_ZNKSt8numpunctIcE9falsenameEv .pdata$_ZNKSt8numpunctIcE9falsenameEv .xdata$_ZNSt15numpunct_bynameIcEC2EPKcy .pdata$_ZNSt15numpunct_bynameIcEC2EPKcy .xdata$_ZNSt15numpunct_bynameIcEC1EPKcy .pdata$_ZNSt15numpunct_bynameIcEC1EPKcy .xdata$_Z      NSt15numpunct_bynameIcEC2ERKSsy .pdata$_ZNSt15numpunct_bynameIcEC2ERKSsy .xdata$_ZNSt15numpunct_bynameIcEC1ERKSsy .pdata$_ZNSt15numpunct_bynameIcEC1ERKSsy .xdata$_ZNSt15numpunct_bynameIcED2Ev .pdata$_ZNSt15numpunct_bynameIcED2Ev .xdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11cha      r_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .xdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt7num_putIcSt19ostreambuf_iterat      orIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv .xdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt11__timepunctIcEC2Ey .pdata$_ZNSt11__timepunctIcEC2Ey .xdata$_ZNSt11__timepunctIcEC1Ey .pdata$_ZNSt      11__timepunctIcEC1Ey .xdata$_ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEy .pdata$_ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEy .xdata$_ZNSt11__timepunctIcEC1EPSt17__timepunct_cacheIcEy .pdata$_ZNSt11__timepunctIcEC1EPSt17__timepunct_cacheIcEy .xdata$_ZNSt11__timepunctIcEC2EPiPKcy .pdata$_ZNSt11__timepunctIcEC2EPiPKcy .xdata$_ZNSt11__timepunctIcEC1EPiPKcy .pdata$_ZNSt11__timepunctIcEC1EPiPKcy .xdata$_ZNKSt11__timepunctIcE15_M_date_formatsEPPKc .pdata$_ZNKSt11__timepunctIcE15_M_date_formatsEPPKc .xdata$_ZNKSt11__timepunctIcE15_M_time_formatsEPPKc .pdata$_ZNKSt11__timepunctIcE15_M_time_formatsEPPKc .xdata$_ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc .pdata$_ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc .xdata$_ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc .pdata$_ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc .xdata$_ZNKSt11__timepunctIcE8_M_am_pmEPPKc .pdata$_ZNKSt11__timepunctIcE8_M_am_pmEPPKc .xdata$_ZNKSt11__timepunctIcE7_M_daysEPPKc .pdata$_ZNKSt11__timepunctIcE7_M_daysEPPKc .xdata$_ZNKSt      11__timepunctIcE19_M_days_abbreviatedEPPKc .pdata$_ZNKSt11__timepunctIcE19_M_days_abbreviatedEPPKc .xdata$_ZNKSt11__timepunctIcE9_M_monthsEPPKc .pdata$_ZNKSt11__timepunctIcE9_M_monthsEPPKc .xdata$_ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc .pdata$_ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc .xdata$_ZNSt11__timepunctIcED2Ev .pdata$_ZNSt11__timepunctIcED2Ev .xdata$_ZNSt17__timepunct_cacheIcEC2Ey .pdata$_ZNSt17__timepunct_cacheIcEC2Ey .xdata$_ZNSt17__timepunct_cacheIcEC1Ey .pdata$_ZNSt17__timepunct_cacheIcEC1Ey .xdata$_ZNSt17__timepunct_cacheIcED2Ev .pdata$_ZNSt17__timepunct_cacheIcED2Ev .xdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc .pdata$_ZNKSt8time_pu      tIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc .xdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .pdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .xdata$_ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt15time_put_bynameIcSt19o      streambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .pdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Ey .xdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .pdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Ey .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istream      buf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcy .xd      ata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcy .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2ERKSsy .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1ERKSsy .xdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .pdata$_ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev .xdata$_ZNSt8messagesIcEC2Ey .pdata$_ZNSt8messagesIcEC2Ey .xdata$_ZNSt8messagesIcEC1Ey .pdata$_ZNSt8messagesIcEC1Ey .xdata$_ZNSt8messagesIcEC2EPiPKcy .pdata$_ZNSt8messagesIcEC2EPiPKcy .xdata$_ZNSt8messagesIcEC1EPiPKcy .pdata$_ZNSt8messagesIcEC1EPiPKcy .xdata$_ZNKSt8messagesIcE4openERKSsRKSt6locale .pdata$_ZNKSt8messagesIcE4openERKSsRKSt6locale .xd      ata$_ZNKSt8messagesIcE4openERKSsRKSt6localePKc .pdata$_ZNKSt8messagesIcE4openERKSsRKSt6localePKc .xdata$_ZNKSt8messagesIcE3getEiiiRKSs .pdata$_ZNKSt8messagesIcE3getEiiiRKSs .xdata$_ZNKSt8messagesIcE5closeEi .pdata$_ZNKSt8messagesIcE5closeEi .xdata$_ZNSt8messagesIcED2Ev .pdata$_ZNSt8messagesIcED2Ev .xdata$_ZNKSt8messagesIcE18_M_convert_to_charERKSs .pdata$_ZNKSt8messagesIcE18_M_convert_to_charERKSs .xdata$_ZNKSt8messagesIcE20_M_convert_from_charEPc .pdata$_ZNKSt8messagesIcE20_M_convert_from_charEPc .xdata$_ZNSt15messages_bynameIcEC2EPKcy .pdata$_ZNSt15messages_bynameIcEC2EPKcy .xdata$_ZNSt15messages_bynameIcEC1EPKcy .pdata$_ZNSt15messages_bynameIcEC1EPKcy .xdata$_ZNSt15messages_bynameIcEC2ERKSsy .pdata$_ZNSt15messages_bynameIcEC2ERKSsy .xdata$_ZNSt15messages_bynameIcEC1ERKSsy .pdata$_ZNSt15messages_bynameIcEC1ERKSsy .xdata$_ZNSt15messages_bynameIcED2Ev .pdata$_ZNSt15messages_bynameIcED2Ev .text$_ZNSt12ctype_bynameIcEC2ERKSsy .xdata$_ZNSt12ctype_bynameIcEC2ERKSsy .pdata$_ZNSt12ctype_bynameIcEC2ERKSsy .x      data$_ZNSt14codecvt_bynameIcciEC2EPKcy .pdata$_ZNSt14codecvt_bynameIcciEC2EPKcy .xdata$_ZNSt14codecvt_bynameIcciEC1EPKcy .pdata$_ZNSt14codecvt_bynameIcciEC1EPKcy .xdata$_ZNSt14codecvt_bynameIcciEC2ERKSsy .pdata$_ZNSt14codecvt_bynameIcciEC2ERKSsy .xdata$_ZNSt14codecvt_bynameIcciEC1ERKSsy .pdata$_ZNSt14codecvt_bynameIcciEC1ERKSsy .xdata$_ZNSt14codecvt_bynameIcciED2Ev .pdata$_ZNSt14codecvt_bynameIcciED2Ev .xdata$_ZNSt7collateIcEC2Ey .pdata$_ZNSt7collateIcEC2Ey .xdata$_ZNSt7collateIcEC1Ey .pdata$_ZNSt7collateIcEC1Ey .xdata$_ZNSt7collateIcEC2EPiy .pdata$_ZNSt7collateIcEC2EPiy .xdata$_ZNSt7collateIcEC1EPiy .pdata$_ZNSt7collateIcEC1EPiy .xdata$_ZNKSt7collateIcE7compareEPKcS2_S2_S2_ .pdata$_ZNKSt7collateIcE7compareEPKcS2_S2_S2_ .xdata$_ZNKSt7collateIcE9transformEPKcS2_ .pdata$_ZNKSt7collateIcE9transformEPKcS2_ .xdata$_ZNKSt7collateIcE4hashEPKcS2_ .pdata$_ZNKSt7collateIcE4hashEPKcS2_ .xdata$_ZNSt7collateIcED2Ev .pdata$_ZNSt7collateIcED2Ev .xdata$_ZNSt14collate_bynameIcEC2EPKcy .pdata$_ZNSt14collate_bynameIcEC2      EPKcy .xdata$_ZNSt14collate_bynameIcEC1EPKcy .pdata$_ZNSt14collate_bynameIcEC1EPKcy .xdata$_ZNSt14collate_bynameIcEC2ERKSsy .pdata$_ZNSt14collate_bynameIcEC2ERKSsy .xdata$_ZNSt14collate_bynameIcEC1ERKSsy .pdata$_ZNSt14collate_bynameIcEC1ERKSsy .xdata$_ZNSt14collate_bynameIcED2Ev .pdata$_ZNSt14collate_bynameIcED2Ev .xdata$_ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale .pdata$_ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale .xdata$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ .pdata$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_      getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZSt9use_facetISt7codecvtIcciEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7codecvtIcciEERKT_RKSt6locale .xdata$_ZSt9use_facetISt7collateIcEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7collateIcEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale .xdata$_ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale .pdata$_ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale .xdata$_ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt10moneypunctIcLb1EEERKT_RKSt6locale .pdata$_ZSt9use_facetISt10moneypunctIcLb       1EEERKT_RKSt6locale .xdata$_ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale .pdata$_ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale .xdata$_ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale .pdata$_ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale .xdata$_ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale .pdata$_ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale .xdata$_ZSt9use_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale .pdata$_ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale .xdata$_ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc .pdata$_ZNKSt8time_putIcS!      t19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc .xdata$_ZSt9use_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8messagesIcEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8messagesIcEERKT_RKSt6locale .xdata$_ZSt9has_facetISt5ctypeIcEEbRKSt6locale .pdata$_ZSt9has_facetISt5ctypeIcEEbRKSt6locale .xdata$_ZSt9has_facetISt7codecvtIcciEEbRKSt6locale .pdata$_ZSt9has_facetISt7codecvtIcciEEbRKSt6locale .xdata$_ZSt9has_facetISt7collateIcEEbRKSt6locale .pdata$_ZSt9has_facetISt7collateIcEEbRKSt6locale .xdata$_ZSt9has_facetISt8numpunctIcEEbRKSt6locale .pdata$_ZSt9has_facetISt8numpunctIcEEbRKSt6locale .xdata$_ZSt9has_facetISt7num_putIcSt19ostreambuf_ite"      ratorIcSt11char_traitsIcEEEEbRKSt6locale .pdata$_ZSt9has_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .pdata$_ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale .pdata$_ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale .xdata$_ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .pdata$_ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .pdata$_ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt11__timepunctIcEEbRKSt6locale .pdata$_ZSt9has_facetISt11__timepunctIcEEbRKSt6locale .xdata$_ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale #      .pdata$_ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .pdata$_ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale .xdata$_ZSt9has_facetISt8messagesIcEEbRKSt6locale .pdata$_ZSt9has_facetISt8messagesIcEEbRKSt6locale .xdata$_ZSt14__add_groupingIcEPT_S1_S0_PKcyPKS0_S5_ .pdata$_ZSt14__add_groupingIcEPT_S1_S0_PKcyPKS0_S5_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcycS6_PcS7_Ri .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcycS6_PcS7_Ri .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcycRSt8ios_basePcS9_Ri .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcycRSt8ios_basePcS9_Ri .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs .$      pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs .pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece .pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece .xdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs .pdata$_ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs .xdata$_ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcxx .pdata$_ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcxx .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6_M_padEcxRSt8ios_basePcPKcRi .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char%      _traitsIcEEE6_M_padEcxRSt8ios_basePcPKcRi .xdata$_ZSt13__int_to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .pdata$_ZSt13__int_to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .xdata$_ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .pdata$_ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .xdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale .xdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl .xdata$_ZNKSt7num_putIcSt19ostreambu&      f_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecl .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecl .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_R'      St8ios_basecT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_RSt8ios_basecT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv .pdata$_ZNKSt7num_pu(      tIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ .pdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ .xdata$_ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece .pdata$_ZNKSt7num_putIcSt19o)      streambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istr*      eambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt8time_getIcSt19istreambu+      f_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_Iost,      ateRe .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_-      getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_ge.      tIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_/      RSt8ios_baseRSt12_Ios_IostateRm .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt110      char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .xdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .pdata$_ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateR1      Ss .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSC_ .pdata$_ZNKSt8time_getIcSt19is2      treambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKcSC_ .text.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKSsy .xdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKSsy .pdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIcEC2ERKSsy .text$_ZNSoD1Ev _ZNSoD1Ev .rdata$_ZTVSo .text$_ZNSoD0Ev _ZNSoD0Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEED1Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEED1Ev .rdata$_ZTVSt13basic_ostreamIwSt11char_traitsIwEE .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEED0Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEED0Ev .text$_ZTv0_n24_NSoD1Ev _ZTv0_n24_NSoD1Ev .text$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED1Ev _ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED1Ev .text$_ZTv0_n24_NSoD0Ev _ZTv0_n24_NSoD0Ev .text$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED0Ev _ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED0Ev .text$_ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSoC1E3      PSt15basic_streambufIcSt11char_traitsIcEE _ZNSoC1EPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSoD2Ev _ZNSoD2Ev .text$_ZNSolsEPFRSoS_E _ZNSolsEPFRSoS_E .text$_ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E _ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .text$_ZNSolsEPFRSt8ios_baseS0_E _ZNSolsEPFRSt8ios_baseS0_E .text$_ZNSo8_M_writeEPKcx _ZNSo8_M_writeEPKcx .text$_ZNSo5flushEv _ZNSo5flushEv .text$_ZNSo5tellpEv _ZNSo5tellpEv .text$_ZNSo5seekpESt4fposIiE _ZNSo5seekpESt4fposIiE .text$_ZNSo5seekpExSt12_Ios_Seekdir _ZNSo5seekpExSt12_Ios_Seekdir .text$_ZNSoC2Ev _ZNSoC2Ev .text$_ZNSoC1Ev _ZNSoC1Ev .text$_ZNSoC2ERSd _ZNSoC2ERSd .text$_ZNSoC1ERSd _ZNSoC1ERSd .text$_ZNSoC2EOSo _ZNSoC2EOSo .text$_ZNSoC1EOSo _ZNSoC1EOSo .text$_ZNSoaSEOSo _ZNSoaSEOSo .text$_ZNSo4swapERSo _ZNSo4swapERSo .text$_ZNSo6sentryC2ERSo _ZNSo6sentryC2ERSo .text$_ZNSo6sentryC1ERSo _ZNSo6sentryC1ERSo .text$_ZNSo6sentryD2Ev _ZNSo6sentryD2Ev .text$_ZNSo6sentryD1Ev _ZNSo6sentryD1Ev .text$_ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE 4      _ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSo3putEc _ZNSo3putEc .text$_ZNSo5writeEPKcx _ZNSo5writeEPKcx .text$_ZNKSo6sentrycvbEv _ZNKSo6sentrycvbEv .text$_ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .text$_ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .text$_ZSt5flushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZSt5flushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .text$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .text$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .text$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags .text$_ZStlsIcSt11char_t5      raitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .text$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .text$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw .text$_ZSt16__ostream_insertIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_x _ZSt16__ostream_insertIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_x .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKc _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_6      ES5_PKc .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa .text$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh .text$_ZNSo9_M_insertIlEERSoT_ _ZNSo9_M_insertIlEERSoT_ .text$_ZNSolsEl _ZNSolsEl .text$_ZNSolsEs _ZNSolsEs .text$_ZNSolsEi _ZNSolsEi .text$_ZNSo9_M_insertImEERSoT_ _ZNSo9_M_insertImEERSoT_ .text$_ZNSolsEm _ZNSolsEm .text$_ZNSolsEt _ZNSolsEt .text$_ZNSolsEj _ZNSolsEj .text$_ZNSo9_M_insertIbEERSoT_ _ZNSo9_M_insertIbEERSoT_ .text$_ZNSolsEb _ZNSolsEb .text$_ZNSo9_M_insertIxEERSoT_ _ZNSo9_M_insertIxEERSoT_ .text$_ZNSolsEx _ZNSolsEx .text$_ZNSo9_M_insertIyEERSoT_ _ZNSo9_M_insertIyEERSoT_ .text$_ZNSolsEy _ZNSolsEy .text$_ZNSo9_M_insertIdEERSoT_ _ZNSo9_M_insertIdEERSoT_ .text$_ZNSolsEd _ZNSolsEd .text$_ZNSolsEf _ZNSolsEf .text$_ZNSo9_M_insertIeEERSoT_ _ZNSo9_M_insertIeEERSoT_ .text$_ZNSolsEe _ZNSolsEe .text$_ZNSo9_M_insertIPKvEERSoT_ _ZNSo9_M_insertIPKvEERSoT_ .text$_Z7      NSolsEPKv _ZNSolsEPKv .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E _ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E _ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEED2Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEED2Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRS2_S3_E _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRS2_S3_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt9basic_iosIwS1_ES5_E _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt9basic_iosIwS1_ES5_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt8ios_baseS4_E _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt8ios_baseS4_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE8_M_writeEPKwx _ZNSt13basic_ostreamIwSt11char_traitsIwEE8_M_writeEPKwx .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5flushEv _ZNSt13basic_ostreamIwSt11char_t8      raitsIwEE5flushEv .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5tellpEv _ZNSt13basic_ostreamIwSt11char_traitsIwEE5tellpEv .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpESt4fposIiE _ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpESt4fposIiE .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpExSt12_Ios_Seekdir _ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpExSt12_Ios_Seekdir .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEEC2Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEEC1Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2ERSt14basic_iostreamIwS1_E _ZNSt13basic_ostreamIwSt11char_traitsIwEEC2ERSt14basic_iostreamIwS1_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1ERSt14basic_iostreamIwS1_E _ZNSt13basic_ostreamIwSt11char_traitsIwEEC1ERSt14basic_iostreamIwS1_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EOS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EOS2_ .text$_ZNSt13basic_ostreamIwSt11char_t9      raitsIwEEC1EOS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EOS2_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEEaSEOS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEEaSEOS2_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE4swapERS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE4swapERS2_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC2ERS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC2ERS2_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC1ERS2_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC1ERS2_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD2Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD2Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD1Ev _ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD1Ev .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPSt15basic_streambufIwS1_E _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPSt15basic_streambufIwS1_E .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE3putEw _ZNSt13basic_ostreamIwSt11char_traitsIwEE3putEw .text$_ZNSt13basic_ostream:      IwSt11char_traitsIwEE5writeEPKwx _ZNSt13basic_ostreamIwSt11char_traitsIwEE5writeEPKwx .text$_ZNKSt13basic_ostreamIwSt11char_traitsIwEE6sentrycvbEv _ZNKSt13basic_ostreamIwSt11char_traitsIwEE6sentrycvbEv .text$_ZSt4endlIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ _ZSt4endlIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .text$_ZSt4endsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ _ZSt4endsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .text$_ZSt5flushIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ _ZSt5flushIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St14_;      Resetiosflags .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_Setbase _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St5_Setw _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St5_Setw .text$_ZSt16__ostream_insertIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_x _ZSt16__ostream_insertIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_x .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_S3_ _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_S3_ .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_ _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_ .text$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_c _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_c .text$_ZStlsIwSt11char_traitsIwEERSt13basi<      c_ostreamIT_T0_ES6_PKc _ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKc .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIlEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIlEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEl _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEl .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEs _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEs .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEi _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEi .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertImEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertImEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEm _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEm .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEt _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEt .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEj _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEj .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIbEERS2_T_ _ZNSt13basic_ostre=      amIwSt11char_traitsIwEE9_M_insertIbEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEb _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEb .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIxEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIxEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEx _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEx .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIyEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIyEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEy _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEy .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIdEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIdEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEd _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEd .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEf _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEf .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIeEERS2_T_ _ZNSt13basic_ostreamIwSt>      11char_traitsIwEE9_M_insertIeEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEe _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEe .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIPKvEERS2_T_ _ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIPKvEERS2_T_ .text$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPKv _ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPKv .rdata$_ZTSSo .rdata$_ZTISo .rdata$_ZTSSt13basic_ostreamIwSt11char_traitsIwEE .rdata$_ZTISt13basic_ostreamIwSt11char_traitsIwEE .rdata$_ZTTSo .rdata$_ZTTSt13basic_ostreamIwSt11char_traitsIwEE .xdata$_ZNSoD1Ev .pdata$_ZNSoD1Ev .xdata$_ZNSoD0Ev .pdata$_ZNSoD0Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED1Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED1Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED0Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED0Ev .xdata$_ZTv0_n24_NSoD1Ev .pdata$_ZTv0_n24_NSoD1Ev .xdata$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED1Ev .pdata$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED1Ev ?      .xdata$_ZTv0_n24_NSoD0Ev .pdata$_ZTv0_n24_NSoD0Ev .xdata$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED0Ev .pdata$_ZTv0_n24_NSt13basic_ostreamIwSt11char_traitsIwEED0Ev .xdata$_ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSoC1EPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSoC1EPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSoD2Ev .pdata$_ZNSoD2Ev .xdata$_ZNSolsEPFRSoS_E .pdata$_ZNSolsEPFRSoS_E .xdata$_ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .pdata$_ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E .xdata$_ZNSolsEPFRSt8ios_baseS0_E .pdata$_ZNSolsEPFRSt8ios_baseS0_E .xdata$_ZNSo8_M_writeEPKcx .pdata$_ZNSo8_M_writeEPKcx .xdata$_ZNSo5flushEv .pdata$_ZNSo5flushEv .xdata$_ZNSo5tellpEv .pdata$_ZNSo5tellpEv .xdata$_ZNSo5seekpESt4fposIiE .pdata$_ZNSo5seekpESt4fposIiE .xdata$_ZNSo5seekpExSt12_Ios_Seekdir .pdata$_ZNSo5seekpExSt12_Ios_Seekdir .xdata$_ZNSoC2Ev .pdata$_ZNSoC2Ev .xdata$_ZNSoC1Ev .pdata$_ZNSoC1Ev .xdata$_ZNSoC2@      ERSd .pdata$_ZNSoC2ERSd .xdata$_ZNSoC1ERSd .pdata$_ZNSoC1ERSd .xdata$_ZNSoC2EOSo .pdata$_ZNSoC2EOSo .xdata$_ZNSoC1EOSo .pdata$_ZNSoC1EOSo .xdata$_ZNSoaSEOSo .pdata$_ZNSoaSEOSo .xdata$_ZNSo4swapERSo .pdata$_ZNSo4swapERSo .xdata$_ZNSo6sentryC2ERSo .pdata$_ZNSo6sentryC2ERSo .xdata$_ZNSo6sentryC1ERSo .pdata$_ZNSo6sentryC1ERSo .xdata$_ZNSo6sentryD2Ev .pdata$_ZNSo6sentryD2Ev .xdata$_ZNSo6sentryD1Ev .pdata$_ZNSo6sentryD1Ev .xdata$_ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE .pdata$_ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE .xdata$_ZNSo3putEc .pdata$_ZNSo3putEc .xdata$_ZNSo5writeEPKcx .pdata$_ZNSo5writeEPKcx .xdata$_ZNKSo6sentrycvbEv .pdata$_ZNKSo6sentrycvbEv .xdata$_ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZSt5flushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt5fA      lushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .xdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw .pdata$_ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw .xdata$_ZSt16__ostream_insertIcSt1B      1char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_x .pdata$_ZSt16__ostream_insertIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_x .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKc .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKc .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa .xdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh .pdata$_ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh .xdata$_ZNSo9_M_insertIlEERSoT_ .pdata$_ZNSo9_M_insertIlEERSoT_ .xdata$_ZNSolsEl .pdata$_ZNSolsEl .xdata$_ZNSolsEs .pdata$_ZNSolsEs .xdaC      ta$_ZNSolsEi .pdata$_ZNSolsEi .xdata$_ZNSo9_M_insertImEERSoT_ .pdata$_ZNSo9_M_insertImEERSoT_ .xdata$_ZNSolsEm .pdata$_ZNSolsEm .xdata$_ZNSolsEt .pdata$_ZNSolsEt .xdata$_ZNSolsEj .pdata$_ZNSolsEj .xdata$_ZNSo9_M_insertIbEERSoT_ .pdata$_ZNSo9_M_insertIbEERSoT_ .xdata$_ZNSolsEb .pdata$_ZNSolsEb .xdata$_ZNSo9_M_insertIxEERSoT_ .pdata$_ZNSo9_M_insertIxEERSoT_ .xdata$_ZNSolsEx .pdata$_ZNSolsEx .xdata$_ZNSo9_M_insertIyEERSoT_ .pdata$_ZNSo9_M_insertIyEERSoT_ .xdata$_ZNSolsEy .pdata$_ZNSolsEy .xdata$_ZNSo9_M_insertIdEERSoT_ .pdata$_ZNSo9_M_insertIdEERSoT_ .xdata$_ZNSolsEd .pdata$_ZNSolsEd .xdata$_ZNSolsEf .pdata$_ZNSolsEf .xdata$_ZNSo9_M_insertIeEERSoT_ .pdata$_ZNSo9_M_insertIeEERSoT_ .xdata$_ZNSolsEe .pdata$_ZNSolsEe .xdata$_ZNSo9_M_insertIPKvEERSoT_ .pdata$_ZNSo9_M_insertIPKvEERSoT_ .xdata$_ZNSolsEPKv .pdata$_ZNSolsEPKv .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EPSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_ostreamIwSt11cD      har_traitsIwEEC1EPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EPSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED2Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEED2Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRS2_S3_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRS2_S3_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt9basic_iosIwS1_ES5_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt9basic_iosIwS1_ES5_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt8ios_baseS4_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPFRSt8ios_baseS4_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE8_M_writeEPKwx .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE8_M_writeEPKwx .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5flushEv .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5flushEv .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5tellpEv .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5tellpEv .xdata$_ZNSt13baE      sic_ostreamIwSt11char_traitsIwEE5seekpESt4fposIiE .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpESt4fposIiE .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpExSt12_Ios_Seekdir .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5seekpExSt12_Ios_Seekdir .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2ERSt14basic_iostreamIwS1_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2ERSt14basic_iostreamIwS1_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1ERSt14basic_iostreamIwS1_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1ERSt14basic_iostreamIwS1_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EOS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC2EOS2_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EOS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEC1EOS2_ .xdata$_ZNF      St13basic_ostreamIwSt11char_traitsIwEEaSEOS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEEaSEOS2_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC2ERS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC2ERS2_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC1ERS2_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryC1ERS2_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD2Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD2Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD1Ev .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE6sentryD1Ev .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPSt15basic_streambufIwS1_E .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPSt15basic_streambufIwS1_E .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE3putEw .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE3putEw .xdata$_ZNSt13basic_ostreamIwSt11char_G      traitsIwEE5writeEPKwx .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE5writeEPKwx .xdata$_ZNKSt13basic_ostreamIwSt11char_traitsIwEE6sentrycvbEv .pdata$_ZNKSt13basic_ostreamIwSt11char_traitsIwEE6sentrycvbEv .xdata$_ZSt4endlIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt4endlIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZSt4endsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt4endsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZSt5flushIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .pdata$_ZSt5flushIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_ .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags .pdata$_ZStlsIwH      St11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St8_Setbase .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St5_Setw .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_St5_Setw .xdata$_ZSt16__ostream_insertIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_x .pdata$_ZSt16__ostream_insertIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_x .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_S3_ .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_S3_ .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_ .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKS3_ .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_I      c .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_c .xdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKc .pdata$_ZStlsIwSt11char_traitsIwEERSt13basic_ostreamIT_T0_ES6_PKc .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIlEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIlEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEl .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEl .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEs .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEs .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEi .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEi .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertImEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertImEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEm .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEm .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEt .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEt .xdata$_ZNStJ      13basic_ostreamIwSt11char_traitsIwEElsEj .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEj .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIbEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIbEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEb .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEb .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIxEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIxEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEx .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEx .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIyEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIyEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEy .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEy .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIdEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIdEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEdK       .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEd .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEf .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEf .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIeEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIeEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEe .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEe .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIPKvEERS2_T_ .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEE9_M_insertIPKvEERS2_T_ .xdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPKv .pdata$_ZNSt13basic_ostreamIwSt11char_traitsIwEElsEPKv _ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ _ZN9__gnu_cxx15__concat_size_tEPcyy _ZN9__gnu_cxx15__snprintf_liteEPcyPKcS0_ .text$_ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ .xdata$_ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ .pdata$_ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ .text$_ZN9__gnu_cxx15__concat_size_tEPcyy .xdata$_ZN9__gnu_cxx15__cL      oncat_size_tEPcyy .pdata$_ZN9__gnu_cxx15__concat_size_tEPcyy .text$_ZN9__gnu_cxx15__snprintf_liteEPcyPKcS0_ .xdata$_ZN9__gnu_cxx15__snprintf_liteEPcyPKcS0_ .pdata$_ZN9__gnu_cxx15__snprintf_liteEPcyPKcS0_ .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcx _ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE4syncEv _ZNSt15basic_streambufIcSt11char_traitsIcEE4syncEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE9showmanycEv _ZNSt15basic_streambufIcSt11char_traitsIcEE9showmaM      nycEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv _ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi _ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi _ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5imbueERKSt6locale _ZNSt15basic_streambufIwSt11char_traitsIwEE5imbueERKSt6locale .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6setbufEPwx _ZNSt15basic_streambufIwSt11char_traitsIwEE6setbufEPwx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt15basic_streambufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode _ZNSt15basic_streambufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE4syncEv _ZNSt15baN      sic_streambufIwSt11char_traitsIwEE4syncEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE9showmanycEv _ZNSt15basic_streambufIwSt11char_traitsIwEE9showmanycEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE9underflowEv _ZNSt15basic_streambufIwSt11char_traitsIwEE9underflowEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pbackfailEt _ZNSt15basic_streambufIwSt11char_traitsIwEE9pbackfailEt .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE8overflowEt _ZNSt15basic_streambufIwSt11char_traitsIwEE8overflowEt .text$_ZNSt15basic_streambufIcSt11char_traitsIcEED1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEED1Ev .rdata$_ZTVSt15basic_streambufIcSt11char_traitsIcEE .text$_ZNSt15basic_streambufIwSt11char_traitsIwEED1Ev _ZNSt15basic_streambufIwSt11char_traitsIwEED1Ev .rdata$_ZTVSt15basic_streambufIwSt11char_traitsIwEE .text$_ZNSt15basic_streambufIcSt11char_traitsIcEED0Ev _ZNSt15basic_streambufIcSt11char_traitsIcEED0Ev .text$_ZNSt15basic_streambufIwSt11char_traitsIwEED0Ev _ZNSt15basic_streambufIwSt11char_traitsIO      wEED0Ev .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcx _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsputnEPKwx _ZNSt15basic_streambufIwSt11char_traitsIwEE6xsputnEPKwx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5uflowEv _ZNSt15basic_streambufIwSt11char_traitsIwEE5uflowEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv _ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcx _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsgetnEPwx _ZNSt15basic_streambufIwSt11char_traitsIwEE6xsgetnEPwx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEED2Ev _ZNSt15basic_streambufIcSt11char_traitsIcEED2Ev .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale _ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE6getlocEv _ZNKSt15basic_streambuP      fIcSt11char_traitsIcEE6getlocEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcx _ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposIiESt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv _ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE8in_availEv _ZNSt15basic_streambufIcSt11char_traitsIcEE8in_availEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv _ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv _ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv .text$_ZNSt15basic_streambufIcSt11char_traitsIQ      cEE5sgetcEv _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetcEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcx _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc _ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv _ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcx _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEEC2Ev _ZNSt15basic_streambufIcSt11char_traitsIcEEC2Ev .text$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEEC1Ev .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE4gptrEv _ZNKStR      15basic_streambufIcSt11char_traitsIcEE4gptrEv .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi _ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ _ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE4pptrEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE4pptrEv .text$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi _ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ _ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE6stosscEv _ZNSt15S      basic_streambufIcSt11char_traitsIcEE6stosscEv .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEx _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEx _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEx .text$_ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ .text$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1ERKS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEEC1ERKS2_ .text$_ZNSt15basic_streambufIcSt11char_traitsIcEEaSERKS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEEaSERKS2_ .text$_ZNSt15basic_streambufIcSt11char_traitsIcEE4swapERS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEE4swapERS2_ .text$_ZSt17__copy_streambufsIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_ _ZSt17__copy_streambufsIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_ .text$_ZNSt15basic_streambufIwSt11char_traitsIwEED2Ev _ZNSt15basic_streambufIwSt11char_traitsIwEED2Ev .text$_ZNSt15bT      asic_streambufIwSt11char_traitsIwEE8pubimbueERKSt6locale _ZNSt15basic_streambufIwSt11char_traitsIwEE8pubimbueERKSt6locale .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE6getlocEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE6getlocEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pubsetbufEPwx _ZNSt15basic_streambufIwSt11char_traitsIwEE9pubsetbufEPwx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekposESt4fposIiESt13_Ios_Openmode _ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekposESt4fposIiESt13_Ios_Openmode .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE7pubsyncEv _ZNSt15basic_streambufIwSt11char_traitsIwEE7pubsyncEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE8in_availEv _ZNSt15basic_streambufIwSt11char_traitsIwEE8in_availEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6snextcEv _ZNSt15U      basic_streambufIwSt11char_traitsIwEE6snextcEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6sbumpcEv _ZNSt15basic_streambufIwSt11char_traitsIwEE6sbumpcEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetcEv _ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetcEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetnEPwx _ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetnEPwx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE9sputbackcEw _ZNSt15basic_streambufIwSt11char_traitsIwEE9sputbackcEw .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE7sungetcEv _ZNSt15basic_streambufIwSt11char_traitsIwEE7sungetcEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputcEw _ZNSt15basic_streambufIwSt11char_traitsIwEE5sputcEw .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputnEPKwx _ZNSt15basic_streambufIwSt11char_traitsIwEE5sputnEPKwx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2Ev _ZNSt15basic_streambufIwSt11char_traitsIwEEC2Ev .text$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1Ev _ZNSt15basic_streambV      ufIwSt11char_traitsIwEEC1Ev .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5ebackEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE5ebackEv .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4gptrEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE4gptrEv .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5egptrEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE5egptrEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5gbumpEi _ZNSt15basic_streambufIwSt11char_traitsIwEE5gbumpEi .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setgEPwS3_S3_ _ZNSt15basic_streambufIwSt11char_traitsIwEE4setgEPwS3_S3_ .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5pbaseEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE5pbaseEv .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4pptrEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE4pptrEv .text$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5epptrEv _ZNKSt15basic_streambufIwSt11char_traitsIwEE5epptrEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE5pbumpEi _ZNSt15basic_streambufIwSt11chW      ar_traitsIwEE5pbumpEi .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setpEPwS3_ _ZNSt15basic_streambufIwSt11char_traitsIwEE4setpEPwS3_ .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE6stosscEv _ZNSt15basic_streambufIwSt11char_traitsIwEE6stosscEv .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_gbumpEx _ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_gbumpEx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_pbumpEx _ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_pbumpEx .text$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2ERKS2_ _ZNSt15basic_streambufIwSt11char_traitsIwEEC2ERKS2_ .text$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1ERKS2_ _ZNSt15basic_streambufIwSt11char_traitsIwEEC1ERKS2_ .text$_ZNSt15basic_streambufIwSt11char_traitsIwEEaSERKS2_ _ZNSt15basic_streambufIwSt11char_traitsIwEEaSERKS2_ .text$_ZNSt15basic_streambufIwSt11char_traitsIwEE4swapERS2_ _ZNSt15basic_streambufIwSt11char_traitsIwEE4swapERS2_ .text$_ZSt17__copy_streambufsIwSt11char_traitsIwEExPSt15basic_streambuX      fIT_T0_ES6_ _ZSt17__copy_streambufsIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_ .rdata$_ZTSSt15basic_streambufIcSt11char_traitsIcEE .rdata$_ZTISt15basic_streambufIcSt11char_traitsIcEE .rdata$_ZTSSt15basic_streambufIwSt11char_traitsIwEE .rdata$_ZTISt15basic_streambufIwSt11char_traitsIwEE .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4syncEv .pdata$_ZNSt15basic_streambufIcSt11chaY      r_traitsIcEE4syncEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9showmanycEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9showmanycEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5imbueERKSt6locale .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5imbueERKSt6locale .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6setbufEPwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6setbufEPwx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIwSt11char_traiZ      tsIwEE7seekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7seekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4syncEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4syncEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9showmanycEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9showmanycEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9underflowEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9underflowEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pbackfailEt .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pbackfailEt .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8overflowEt .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8overflowEt .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEED1Ev .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEED1Ev .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED1Ev .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED1Ev .xdata$_ZNSt15basic_streambufIcSt11char_traitsIc[      EED0Ev .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEED0Ev .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED0Ev .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED0Ev .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsputnEPKwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsputnEPKwx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5uflowEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5uflowEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsgetnEPwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6xsgetnEPwx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEED2Ev .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEED2E\      v .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE6getlocEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE6getlocEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8in_availEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE8in_av]      ailEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetcEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetcEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcx .xdata$_ZNSt15basic_streambufIcSt11char_^      traitsIcEEC2Ev .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC2Ev .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1Ev .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1Ev .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE4gptrEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE4gptrEv .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE4pptrEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE_      4pptrEv .xdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv .pdata$_ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6stosscEv .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE6stosscEv .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEx .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEx .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1ERKS2_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEC1ERKS2_ .xdata$_ZNSt15basic_st`      reambufIcSt11char_traitsIcEEaSERKS2_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEEaSERKS2_ .xdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4swapERS2_ .pdata$_ZNSt15basic_streambufIcSt11char_traitsIcEE4swapERS2_ .xdata$_ZSt17__copy_streambufsIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_ .pdata$_ZSt17__copy_streambufsIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_ .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED2Ev .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEED2Ev .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8pubimbueERKSt6locale .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8pubimbueERKSt6locale .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE6getlocEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE6getlocEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pubsetbufEPwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9pubsetbufEPwx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .pdata$_ZNSt15basic_streambua      fIwSt11char_traitsIwEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekposESt4fposIiESt13_Ios_Openmode .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE10pubseekposESt4fposIiESt13_Ios_Openmode .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7pubsyncEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7pubsyncEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8in_availEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE8in_availEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6snextcEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6snextcEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6sbumpcEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6sbumpcEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetcEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetcEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetnEPwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sgetnEPwx .xdata$_ZNSt15basic_streambufIwSt11chab      r_traitsIwEE9sputbackcEw .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE9sputbackcEw .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7sungetcEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE7sungetcEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputcEw .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputcEw .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputnEPKwx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5sputnEPKwx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2Ev .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2Ev .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1Ev .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1Ev .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5ebackEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5ebackEv .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4gptrEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4gptrEv .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5egptrEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitc      sIwEE5egptrEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5gbumpEi .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5gbumpEi .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setgEPwS3_S3_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setgEPwS3_S3_ .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5pbaseEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5pbaseEv .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4pptrEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE4pptrEv .xdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5epptrEv .pdata$_ZNKSt15basic_streambufIwSt11char_traitsIwEE5epptrEv .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5pbumpEi .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE5pbumpEi .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setpEPwS3_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4setpEPwS3_ .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6stosscEv .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE6stosscEv .xdata$_ZNSt15basic_streambufIwSt1d      1char_traitsIwEE12__safe_gbumpEx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_gbumpEx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_pbumpEx .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE12__safe_pbumpEx .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2ERKS2_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC2ERKS2_ .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1ERKS2_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEC1ERKS2_ .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEaSERKS2_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEEaSERKS2_ .xdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4swapERS2_ .pdata$_ZNSt15basic_streambufIwSt11char_traitsIwEE4swapERS2_ .xdata$_ZSt17__copy_streambufsIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_ .pdata$_ZSt17__copy_streambufsIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc .texe      t$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv .text$_ZNSf      t7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_g      M_get_allocatorEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_S_assignEPcyc _ZNSt7__cxx1112basic_stringIcSt11char_th      raitsIcESaIcEE9_S_assignEPcyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcS4_EESA_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcS4_EESA_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcS5_S5_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcS5_S5_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsi      IcESaIcEE9_M_assignERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_assignERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2Ev _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2Ev .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1Ev _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1Ev .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EycRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EycRKj      S3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EycRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EycRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED2Ev _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED2Ev .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED1Ev _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED1Ev .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSERKS4_ _ZNSt7__cxx1112basic_stringIcSt11ck      har_traitsIcESaIcEEaSERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv _ZNSt7__cxxl      1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv .text$_ZNKSt7__cxx1112basic_stringIcSt11m      char_traitsIcESaIcEE8max_sizeEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8max_sizeEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESn      aIcEEixEy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9push_backEc _ZNSt7__cxx1112basic_stringIcSt11char_traio      tsIcESaIcEE9push_backEc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv .text$_ZNSt7__cxx1112basic_sp      tringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratoq      rIPKcS4_EEc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replaceEyyPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replaceEyyPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy .text$_ZNSt7__cxx1112basic_stringIr      cSt11char_traitsIcESaIcEE6assignEPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ .text$_ZNSt7__cxx1112bs      asic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_t      cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_yy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_yy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7u      replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy _ZNSt7__cxx1112basiv      c_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendESt16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEw      St16initializer_listIcE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5c_strEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5c_strEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy .text$x      _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEy      13find_first_ofEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcyy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12z      find_last_ofEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy .text$_ZNKSt7__cxx1112basi{      c_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEcy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEPKc _ZNKSt7__cxx1112basic_stringIcSt11char_|      traitsIcESaIcEE7compareEPKc .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKcy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcOS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcOS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcOS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcOS3_ .text$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112bas}      ic_stringIT_T0_T1_EEPKS5_RKS8_ _ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .text$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ _ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvT_SA_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvT_SA_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .text$_ZNSt7__cxx1~      112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKcS4_EEEEvT_SB_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKcS4_EEEEvT_SB_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPcEEvT_S7_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPcEEvT_S7_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERK      S4_ .text$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ _ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPcvEET_S7_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPcvEET_S7_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPcvEET_S7_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPcvEET_S7_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPKcEEvT_S8_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPKcEEvT_S8_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcES�      aIcEEC2ERKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yyRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yyRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yyRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yyRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcyRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcyRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcyRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcyRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcRKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcRKS3_ _ZNSt7__cxx1112basic_stringIcSt�      11char_traitsIcESaIcEEC1EPKcRKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ESt16initializer_listIcERKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ESt16initializer_listIcERKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ESt16initializer_listIcERKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ESt16initializer_listIcERKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPKcvEET_S8_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPKcvEET_S8_RKS3_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPKcvEET_S8_RKS3_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPKcvEET_S8_RKS3_ .text$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy _ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy .text$_ZN9__gnu_cxxeqIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ _ZN9__gnu_cxxeqIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRK�      NS_17__normal_iteratorIT_T0_EESD_ .text$_ZN9__gnu_cxxeqIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ _ZN9__gnu_cxxeqIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ .rdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4nposE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEPc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_lengthEy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_M_dataEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .pdata$_ZNKSt7__cxx1�      112basic_stringIcSt11char_traitsIcESaIcEE13_M_local_dataEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_capacityEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_M_set_lengthEy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_is_localEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_createERyy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_disposeEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_destroyEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_�      traitsIcESaIcEE12_M_constructEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE18_M_construct_aux_2Eyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16_M_get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_checkEyPKc .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE15_M_check_lengthEyyPKc .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy .pdata$_ZNKSt7_�      _cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_limitEyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE11_M_disjunctEPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_copyEPcPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7_S_moveEPcPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_S_assignEPcyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_S_assignEPcyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_i�      teratorIPKcS4_EESA_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcS4_EESA_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcS5_S5_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcS5_S5_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13_S_copy_charsEPcPKcS7_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_S_compareEyy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_assignERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_assignERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_mutateEyyPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy �      .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8_M_eraseEyy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2Ev .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2Ev .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1Ev .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1Ev .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EycRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EycRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EycRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EycRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcES�      aIcEEC2EOS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EOS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EOS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED2Ev .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED2Ev .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED1Ev .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEED1Ev .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEOS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11c�      har_traitsIcESaIcEE5beginEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5beginEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE3endEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6rbeginEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4rendEv .pdata$_ZNKSt7__cxx111�      2basic_stringIcSt11char_traitsIcESaIcEE4rendEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6cbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4cendEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7crbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5crendEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4sizeEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6lengthEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8max_sizeEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traits�      IcESaIcEE8max_sizeEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8capacityEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7reserveEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13shrink_to_fitEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5clearEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5emptyEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEixEy .xdata$_ZNK�      St7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE2atEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5frontEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4backEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9push_backEc .pdata�      $_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9push_backEc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEOS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEyy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv .pdata$_Z�      NSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE8pop_backEv .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE14_M_replace_auxEyyyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6resizeEy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc .pdata$_ZNSt7__cxx111�      2basic_stringIcSt11char_traitsIcESaIcEE6insertEyyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_yc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPKcS4_EEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replaceEyyPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE10_M_replac�      eEyyPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSESt16initializer_listIcE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignESt16initializer_listIcE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6assignEPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcES�      aIcEEaSEPKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEaSEPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_RKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_y .xdata$_ZNSt7__cxx1�      112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_PcSA_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_S8_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_St16initializer_listIcE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyRKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyRKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7r�      eplaceEyyRKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_NS6_IPcS4_EESB_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S9_S9_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EESt16initializer_listIcE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEyyPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEyPKc .pdata$_ZNSt7__cxx1112basi�      c_stringIcSt11char_traitsIcESaIcEE6insertEyPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPKcS4_EES9_S8_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE9_M_appendEPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKcy .xd�      ata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendEPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLEPKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendESt16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6appendESt16initializer_listIcE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEpLESt16initializer_listIcE .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4copyEPcyy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4swapERS4_ .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5c_strEv .pdata$_ZNKSt7__cxx1112basi�      c_stringIcSt11char_traitsIcESaIcEE5c_strEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4dataEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEPKcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4findEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy .pdata$_ZNKSt7__cxx1112ba�      sic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEPKcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5rfindEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEPKcy .xdata$_ZNKSt7__cxx1112basic_st�      ringIcSt11char_traitsIcESaIcEE13find_first_ofEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE13find_first_ofEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEPKcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12find_last_ofEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17�      find_first_not_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEPKcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE17find_first_not_ofEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcyy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEPKcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_t�      raitsIcESaIcEE16find_last_not_ofEcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE16find_last_not_ofEcy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareERKS4_ .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_ .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyRKS4_yy .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEPKc .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEPKc .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKc .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7compareEyyPKcy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traits�      IcESaIcEE7compareEyyPKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcOS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC2EPcOS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcOS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_Alloc_hiderC1EPcOS3_ .xdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .pdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .xdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ .pdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_s�      tringIT_T0_T1_EES5_RKS8_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvT_SA_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvT_SA_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IN9__gnu_cxx17__normal_iteratorIPcS4_EEvEET_SA_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKcS4_EEEEvT_SB_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIN9__gnu_cxx17__no�      rmal_iteratorIPKcS4_EEEEvT_SB_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPcEEvT_S7_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPcEEvT_S7_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_ .xdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .pdata$_ZStplIcSt11char_traitsIcESaIcEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .�      xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPcvEET_S7_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPcvEET_S7_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPcvEET_S7_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPcvEET_S7_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPKcEEvT_S8_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE12_M_constructIPKcEEvT_S8_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcS�      t11char_traitsIcESaIcEEC1ERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ERKS4_yyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ERKS4_yyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2EPKcRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1EPKcRKS3_ .xdata$_ZNSt7__cxx1112basic�      _stringIcSt11char_traitsIcESaIcEEC2ESt16initializer_listIcERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2ESt16initializer_listIcERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ESt16initializer_listIcERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1ESt16initializer_listIcERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPKcvEET_S8_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC2IPKcvEET_S8_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPKcvEET_S8_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEC1IPKcvEET_S8_RKS3_ .xdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy .pdata$_ZNKSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6substrEyy .xdata$_ZN9__gnu_cxxeqIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ .pdata$_ZN9__gnu_cxxeqIPcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal�      _iteratorIT_T0_EESD_ .xdata$_ZN9__gnu_cxxeqIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ .pdata$_ZN9__gnu_cxxeqIPKcNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ .text$_ZNKSt10moneypunctIwLb0EE16do_decimal_pointEv _ZNKSt10moneypunctIwLb0EE16do_decimal_pointEv .text$_ZNKSt10moneypunctIwLb0EE16do_thousands_sepEv _ZNKSt10moneypunctIwLb0EE16do_thousands_sepEv .text$_ZNKSt10moneypunctIwLb0EE14do_frac_digitsEv _ZNKSt10moneypunctIwLb0EE14do_frac_digitsEv .text$_ZNKSt10moneypunctIwLb0EE13do_pos_formatEv _ZNKSt10moneypunctIwLb0EE13do_pos_formatEv .text$_ZNKSt10moneypunctIwLb0EE13do_neg_formatEv _ZNKSt10moneypunctIwLb0EE13do_neg_formatEv .text$_ZNKSt10moneypunctIwLb1EE16do_decimal_pointEv _ZNKSt10moneypunctIwLb1EE16do_decimal_pointEv .text$_ZNKSt10moneypunctIwLb1EE16do_thousands_sepEv _ZNKSt10moneypunctIwLb1EE16do_thousands_sepEv .text$_ZNKSt10moneypunctIwLb1EE14do_frac_digitsEv _ZNKSt10moneypunctIwLb1EE14do_frac_digits�      Ev .text$_ZNKSt10moneypunctIwLb1EE13do_pos_formatEv _ZNKSt10moneypunctIwLb1EE13do_pos_formatEv .text$_ZNKSt10moneypunctIwLb1EE13do_neg_formatEv _ZNKSt10moneypunctIwLb1EE13do_neg_formatEv .text$_ZNSt17moneypunct_bynameIwLb0EED1Ev _ZNSt17moneypunct_bynameIwLb0EED1Ev .rdata$_ZTVSt17moneypunct_bynameIwLb0EE .text$_ZNSt17moneypunct_bynameIwLb1EED1Ev _ZNSt17moneypunct_bynameIwLb1EED1Ev .rdata$_ZTVSt17moneypunct_bynameIwLb1EE .text$_ZNKSt8numpunctIwE16do_decimal_pointEv _ZNKSt8numpunctIwE16do_decimal_pointEv .text$_ZNKSt8numpunctIwE16do_thousands_sepEv _ZNKSt8numpunctIwE16do_thousands_sepEv .text$_ZNSt15numpunct_bynameIwED1Ev _ZNSt15numpunct_bynameIwED1Ev .rdata$_ZTVSt15numpunct_bynameIwE .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .text$_ZNKSt8messagesIwE7do_openERKSsRKSt6locale _ZNKSt8messagesIwE7do_openERKSsRKSt6locale .text$_ZNKSt8messagesIwE8do_closeEi _ZNKSt8messagesIwE8do_closeEi .�      text$_ZNKSt7collateIwE7do_hashEPKwS2_ _ZNKSt7collateIwE7do_hashEPKwS2_ .text$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt17__timepunct_cacheIwED1Ev _ZNSt17__timepunct_cacheIwED1Ev .rdata$_ZTVSt17__timepunct_cacheIwE .text$_�      ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .rdata$_ZTVSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .text$_ZNSt17moneypunct_bynameIwLb0EED0Ev _ZNSt17moneypunct_bynameIwLb0EED0Ev .text$_ZNSt17moneypunct_bynameIwLb1EED0Ev _ZNSt17moneypunct_bynameIwLb1EED0Ev .text$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .te�      xt$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt15numpunct_bynameIwED0Ev _ZNSt15numpunct_bynameIwED0Ev .text$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt17__timepunct_cacheIwED0Ev _ZNSt17__timepunct_cacheIwED0Ev .text$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNSt15time_get_bynameIwSt19istream�      buf_iteratorIwSt11char_traitsIwEEED0Ev _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .text$_ZNKSt10moneypunctIwLb0EE11do_groupingEv _ZNKSt10moneypunctIwLb0EE11do_groupingEv .text$_ZNKSt10moneypunctIwLb1EE11do_groupingEv _ZNKSt10moneypunctIwLb1EE11do_groupingEv .text$_ZNKSt8numpunctIwE11do_groupingEv _ZNKSt8numpunctIwE11do_groupingEv .text$_ZNKSt10moneypunctIwLb0EE14do_curr_symbolEv _ZNKSt10moneypunctIwLb0EE14do_curr_symbolEv .text$_ZNKSt10moneypunctIwLb0EE16do_positive_signEv _ZNKSt10moneypunctIwLb0EE16do_positive_signEv .text$_ZNKSt10moneypunctIwLb0EE16do_negative_signEv _ZNKSt10moneypunctIwLb0EE16do_negative_signEv .text$_ZNKSt10moneypunctIwLb1EE14do_curr_symbolEv _ZNKSt10moneypunctIwLb1EE14do_curr_symbolEv .text$_ZNKSt10moneypunctIwLb1EE16do_positive_signEv _ZNKSt10moneypunctIwLb1EE16do_positive_signEv .text$_ZNKSt10moneypunctIwLb1EE16do_negative_signEv _ZNKSt10moneypunctIwLb1EE16do_negative_signEv .text$_ZNKSt8numpunctIwE11do_truenameEv _ZNKSt8numpunctIwE11do_truenameEv�       .text$_ZNKSt8numpunctIwE12do_falsenameEv _ZNKSt8numpunctIwE12do_falsenameEv .text$_ZNSt8messagesIwED1Ev _ZNSt8messagesIwED1Ev .rdata$_ZTVSt8messagesIwE .text$_ZNSt8messagesIwED0Ev _ZNSt8messagesIwED0Ev .text$_ZNSt7collateIwED1Ev _ZNSt7collateIwED1Ev .rdata$_ZTVSt7collateIwE .text$_ZNSt7collateIwED0Ev _ZNSt7collateIwED0Ev .text$_ZNSt15messages_bynameIwED1Ev _ZNSt15messages_bynameIwED1Ev .text$_ZNSt15messages_bynameIwED0Ev _ZNSt15messages_bynameIwED0Ev .text$_ZNSt14collate_bynameIwED1Ev _ZNSt14collate_bynameIwED1Ev .text$_ZNSt14collate_bynameIwED0Ev _ZNSt14collate_bynameIwED0Ev .text$_ZNSt11__timepunctIwED1Ev _ZNSt11__timepunctIwED1Ev .rdata$_ZTVSt11__timepunctIwE .text$_ZNSt11__timepunctIwED0Ev _ZNSt11__timepunctIwED0Ev .text$_ZNSt14codecvt_bynameIwciED1Ev _ZNSt14codecvt_bynameIwciED1Ev .rdata$_ZTVSt14codecvt_bynameIwciE .text$_ZNSt14codecvt_bynameIwciED0Ev _ZNSt14codecvt_bynameIwciED0Ev _ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.43 .text$_ZNKSt7collateIwE12do_transformEPKwS2_ _ZNK�      St7collateIwE12do_transformEPKwS2_ .text$_ZNKSt7collateIwE10do_compareEPKwS2_S2_S2_ _ZNKSt7collateIwE10do_compareEPKwS2_S2_S2_ .text$_ZNSt18__moneypunct_cacheIwLb0EEC2Ey _ZNSt18__moneypunct_cacheIwLb0EEC2Ey .text$_ZNSt18__moneypunct_cacheIwLb0EEC1Ey _ZNSt18__moneypunct_cacheIwLb0EEC1Ey .text$_ZNSt18__moneypunct_cacheIwLb0EED2Ev _ZNSt18__moneypunct_cacheIwLb0EED2Ev .text$_ZNSt18__moneypunct_cacheIwLb1EEC2Ey _ZNSt18__moneypunct_cacheIwLb1EEC2Ey .text$_ZNSt18__moneypunct_cacheIwLb1EEC1Ey _ZNSt18__moneypunct_cacheIwLb1EEC1Ey .text$_ZNSt18__moneypunct_cacheIwLb1EED2Ev _ZNSt18__moneypunct_cacheIwLb1EED2Ev .text$_ZNSt10moneypunctIwLb0EEC2Ey _ZNSt10moneypunctIwLb0EEC2Ey .rdata$_ZTVSt10moneypunctIwLb0EE .text$_ZNSt10moneypunctIwLb0EEC1Ey _ZNSt10moneypunctIwLb0EEC1Ey .text$_ZNSt10moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy _ZNSt10moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .text$_ZNSt10moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy _ZNSt10moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy �      .text$_ZNSt10moneypunctIwLb0EEC2EPiPKcy _ZNSt10moneypunctIwLb0EEC2EPiPKcy .text$_ZNSt10moneypunctIwLb0EEC1EPiPKcy _ZNSt10moneypunctIwLb0EEC1EPiPKcy .text$_ZNKSt10moneypunctIwLb0EE13decimal_pointEv _ZNKSt10moneypunctIwLb0EE13decimal_pointEv .text$_ZNKSt10moneypunctIwLb0EE13thousands_sepEv _ZNKSt10moneypunctIwLb0EE13thousands_sepEv .text$_ZNKSt10moneypunctIwLb0EE8groupingEv _ZNKSt10moneypunctIwLb0EE8groupingEv .text$_ZNKSt10moneypunctIwLb0EE11curr_symbolEv _ZNKSt10moneypunctIwLb0EE11curr_symbolEv .text$_ZNKSt10moneypunctIwLb0EE13positive_signEv _ZNKSt10moneypunctIwLb0EE13positive_signEv .text$_ZNKSt10moneypunctIwLb0EE13negative_signEv _ZNKSt10moneypunctIwLb0EE13negative_signEv .text$_ZNKSt10moneypunctIwLb0EE11frac_digitsEv _ZNKSt10moneypunctIwLb0EE11frac_digitsEv .text$_ZNKSt10moneypunctIwLb0EE10pos_formatEv _ZNKSt10moneypunctIwLb0EE10pos_formatEv .text$_ZNKSt10moneypunctIwLb0EE10neg_formatEv _ZNKSt10moneypunctIwLb0EE10neg_formatEv .text$_ZNSt10moneypunctIwLb1EEC2Ey _ZNSt10moneypunctIwLb1EEC2Ey .rdata$_�      ZTVSt10moneypunctIwLb1EE .text$_ZNSt10moneypunctIwLb1EEC1Ey _ZNSt10moneypunctIwLb1EEC1Ey .text$_ZNSt10moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy _ZNSt10moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .text$_ZNSt10moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy _ZNSt10moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .text$_ZNSt10moneypunctIwLb1EEC2EPiPKcy _ZNSt10moneypunctIwLb1EEC2EPiPKcy .text$_ZNSt10moneypunctIwLb1EEC1EPiPKcy _ZNSt10moneypunctIwLb1EEC1EPiPKcy .text$_ZNKSt10moneypunctIwLb1EE13decimal_pointEv _ZNKSt10moneypunctIwLb1EE13decimal_pointEv .text$_ZNKSt10moneypunctIwLb1EE13thousands_sepEv _ZNKSt10moneypunctIwLb1EE13thousands_sepEv .text$_ZNKSt10moneypunctIwLb1EE8groupingEv _ZNKSt10moneypunctIwLb1EE8groupingEv .text$_ZNKSt10moneypunctIwLb1EE11curr_symbolEv _ZNKSt10moneypunctIwLb1EE11curr_symbolEv .text$_ZNKSt10moneypunctIwLb1EE13positive_signEv _ZNKSt10moneypunctIwLb1EE13positive_signEv .text$_ZNKSt10moneypunctIwLb1EE13negative_signEv _ZNKSt10moneypunctIwLb1EE13negative_si�      gnEv .text$_ZNKSt10moneypunctIwLb1EE11frac_digitsEv _ZNKSt10moneypunctIwLb1EE11frac_digitsEv .text$_ZNKSt10moneypunctIwLb1EE10pos_formatEv _ZNKSt10moneypunctIwLb1EE10pos_formatEv .text$_ZNKSt10moneypunctIwLb1EE10neg_formatEv _ZNKSt10moneypunctIwLb1EE10neg_formatEv .text$_ZNSt17moneypunct_bynameIwLb0EEC2EPKcy _ZNSt17moneypunct_bynameIwLb0EEC2EPKcy .text$_ZNSt17moneypunct_bynameIwLb0EEC1EPKcy _ZNSt17moneypunct_bynameIwLb0EEC1EPKcy .text$_ZNSt17moneypunct_bynameIwLb0EEC2ERKSsy _ZNSt17moneypunct_bynameIwLb0EEC2ERKSsy .text$_ZNSt17moneypunct_bynameIwLb0EEC1ERKSsy _ZNSt17moneypunct_bynameIwLb0EEC1ERKSsy .text$_ZNSt17moneypunct_bynameIwLb0EED2Ev _ZNSt17moneypunct_bynameIwLb0EED2Ev .text$_ZNSt17moneypunct_bynameIwLb1EEC2EPKcy _ZNSt17moneypunct_bynameIwLb1EEC2EPKcy .text$_ZNSt17moneypunct_bynameIwLb1EEC1EPKcy _ZNSt17moneypunct_bynameIwLb1EEC1EPKcy .text$_ZNSt17moneypunct_bynameIwLb1EEC2ERKSsy _ZNSt17moneypunct_bynameIwLb1EEC2ERKSsy .text$_ZNSt17moneypunct_bynameIwLb1EEC1ERKSsy _ZNSt17moneypunct_bynameIwLb1EEC1�      ERKSsy .text$_ZNSt17moneypunct_bynameIwLb1EED2Ev _ZNSt17moneypunct_bynameIwLb1EED2Ev .text$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE .text$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt9money_putIwSt19ostreambuf_iteratorI�      wSt11char_traitsIwEEEC2Ey _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewe _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewe .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewRKSbIwS2_SaIwEE _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .text$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt16__numpunct_cacheIwEC2Ey _ZNSt16__numpunct_cacheIwEC2Ey .text$_ZNSt16__numpunct_cacheIwEC1Ey _ZNSt16__numpunct_cacheIwEC1Ey .text$_ZNSt16__numpunct_cacheIwED2Ev _ZNSt16__numpunct_cacheIwED2Ev .text$_ZNSt8numpunctIwEC2Ey _ZNSt8numpunctIwEC2Ey .�      rdata$_ZTVSt8numpunctIwE .text$_ZNSt8numpunctIwEC1Ey _ZNSt8numpunctIwEC1Ey .text$_ZNSt8numpunctIwEC2EPSt16__numpunct_cacheIwEy _ZNSt8numpunctIwEC2EPSt16__numpunct_cacheIwEy .text$_ZNSt8numpunctIwEC1EPSt16__numpunct_cacheIwEy _ZNSt8numpunctIwEC1EPSt16__numpunct_cacheIwEy .text$_ZNSt8numpunctIwEC2EPiy _ZNSt8numpunctIwEC2EPiy .text$_ZNSt8numpunctIwEC1EPiy _ZNSt8numpunctIwEC1EPiy .text$_ZNKSt8numpunctIwE13decimal_pointEv _ZNKSt8numpunctIwE13decimal_pointEv .text$_ZNKSt8numpunctIwE13thousands_sepEv _ZNKSt8numpunctIwE13thousands_sepEv .text$_ZNKSt8numpunctIwE8groupingEv _ZNKSt8numpunctIwE8groupingEv .text$_ZNKSt8numpunctIwE8truenameEv _ZNKSt8numpunctIwE8truenameEv .text$_ZNKSt8numpunctIwE9falsenameEv _ZNKSt8numpunctIwE9falsenameEv .text$_ZNSt15numpunct_bynameIwEC2EPKcy _ZNSt15numpunct_bynameIwEC2EPKcy .text$_ZNSt15numpunct_bynameIwEC1EPKcy _ZNSt15numpunct_bynameIwEC1EPKcy .text$_ZNSt15numpunct_bynameIwEC2ERKSsy _ZNSt15numpunct_bynameIwEC2ERKSsy .text$_ZNSt15numpunct_bynameIwEC1ERKSsy _ZNSt15numpunct_bynameI�      wEC1ERKSsy .text$_ZNSt15numpunct_bynameIwED2Ev _ZNSt15numpunct_bynameIwED2Ev .text$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .text$_ZNKSt7num_getIwSt1�      9istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .text$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewb _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewb .text$_ZNKSt7num_putIwSt19ost�      reambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewd _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewd .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewe _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewe .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPKv _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPKv .text$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt11__timepunctIwEC2Ey _ZNSt11__timepunctIwEC2Ey .text$_ZNSt11__timepunctIwEC1Ey _ZNSt11__timepunctIwEC1Ey .text$_ZNSt11__timepunctIwEC2EPSt17__timepunct_cacheIwEy _ZNSt11__timepunctIwEC2EPSt17__timepunct_cacheIwEy .text$_ZNSt11__timepunctIwEC1EPSt17__timepunct_cacheIwEy _ZNSt11__timepunctIwEC1EPSt17__timepunct_cacheIwEy .text$_ZNSt11__timepunctIwEC2EPiPKcy _ZNSt11__timep�      unctIwEC2EPiPKcy .text$_ZNSt11__timepunctIwEC1EPiPKcy _ZNSt11__timepunctIwEC1EPiPKcy .text$_ZNKSt11__timepunctIwE15_M_date_formatsEPPKw _ZNKSt11__timepunctIwE15_M_date_formatsEPPKw .text$_ZNKSt11__timepunctIwE15_M_time_formatsEPPKw _ZNKSt11__timepunctIwE15_M_time_formatsEPPKw .text$_ZNKSt11__timepunctIwE20_M_date_time_formatsEPPKw _ZNKSt11__timepunctIwE20_M_date_time_formatsEPPKw .text$_ZNKSt11__timepunctIwE15_M_am_pm_formatEPKw _ZNKSt11__timepunctIwE15_M_am_pm_formatEPKw .text$_ZNKSt11__timepunctIwE8_M_am_pmEPPKw _ZNKSt11__timepunctIwE8_M_am_pmEPPKw .text$_ZNKSt11__timepunctIwE7_M_daysEPPKw _ZNKSt11__timepunctIwE7_M_daysEPPKw .text$_ZNKSt11__timepunctIwE19_M_days_abbreviatedEPPKw _ZNKSt11__timepunctIwE19_M_days_abbreviatedEPPKw .text$_ZNKSt11__timepunctIwE9_M_monthsEPPKw _ZNKSt11__timepunctIwE9_M_monthsEPPKw .text$_ZNKSt11__timepunctIwE21_M_months_abbreviatedEPPKw _ZNKSt11__timepunctIwE21_M_months_abbreviatedEPPKw .text$_ZNSt11__timepunctIwED2Ev _ZNSt11__timepunctIwED2Ev .text$_ZNSt17__timepunct_cach�      eIwEC2Ey _ZNSt17__timepunct_cacheIwEC2Ey .text$_ZNSt17__timepunct_cacheIwEC1Ey _ZNSt17__timepunct_cacheIwEC1Ey .text$_ZNSt17__timepunct_cacheIwED2Ev _ZNSt17__timepunct_cacheIwED2Ev .text$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmcc _ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmcc .text$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .rdata$_ZTVSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsI�      wEEE .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .text$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .text$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv _ZNKSt8time_ge�      tIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8�      time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .rdata$_ZTVSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy _ZNSt15time_get_b�      ynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .text$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev _ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .text$_ZNSt8messagesIwEC2Ey _ZNSt8messagesIwEC2Ey .text$_ZNSt8messagesIwEC1Ey _ZNSt8messagesIwEC1Ey .text$_ZNSt8messagesIwEC2EPiPKcy _ZNSt8messagesIwEC2EPiPKcy .text$_ZNSt8messagesIwEC1EPiPKcy _ZNSt8messagesIwEC1EPiPKcy .text$_ZNKSt8messagesIwE4openERKSsRKSt6locale _ZNKSt8messagesIwE4openERKSsRKSt6locale .text$_ZNKSt8messagesIwE4openERKSsRKSt6localePKc _ZNKSt8messagesIwE4openERKSsRKSt6localePKc .text$_ZNKSt8messagesIwE3getEiiiRKSbIwSt11char_traitsIwESaIwEE _ZNKSt8messagesIwE3getEiiiRKSbIwSt11char_traitsIwESaIwEE .text$_ZNKSt8messagesIwE5closeEi _ZNKSt8messagesIwE5closeEi .text$_ZNSt8messagesIwED2Ev _ZNSt8messagesIwED2Ev .text$_ZNKSt8messagesIwE18_M_convert_to_charERKSbIwSt11char_traitsIwESaIwEE _ZNKSt8messagesIwE18_M_convert_to_charERKSbIwSt11char_traitsIwESaIwEE .text$_ZNKSt8messagesIwE20_�      M_convert_from_charEPc _ZNKSt8messagesIwE20_M_convert_from_charEPc .text$_ZNSt15messages_bynameIwEC2EPKcy _ZNSt15messages_bynameIwEC2EPKcy .rdata$_ZTVSt15messages_bynameIwE .text$_ZNSt15messages_bynameIwEC1EPKcy _ZNSt15messages_bynameIwEC1EPKcy .text$_ZNSt15messages_bynameIwEC2ERKSsy _ZNSt15messages_bynameIwEC2ERKSsy .text$_ZNSt15messages_bynameIwEC1ERKSsy _ZNSt15messages_bynameIwEC1ERKSsy .text$_ZNSt15messages_bynameIwED2Ev _ZNSt15messages_bynameIwED2Ev _ZNSt12ctype_bynameIwEC2ERKSsy _ZNSt12ctype_bynameIwEC1ERKSsy .text$_ZNSt14codecvt_bynameIwciEC2EPKcy _ZNSt14codecvt_bynameIwciEC2EPKcy .text$_ZNSt14codecvt_bynameIwciEC1EPKcy _ZNSt14codecvt_bynameIwciEC1EPKcy .text$_ZNSt14codecvt_bynameIwciEC2ERKSsy _ZNSt14codecvt_bynameIwciEC2ERKSsy .text$_ZNSt14codecvt_bynameIwciEC1ERKSsy _ZNSt14codecvt_bynameIwciEC1ERKSsy .text$_ZNSt14codecvt_bynameIwciED2Ev _ZNSt14codecvt_bynameIwciED2Ev .text$_ZNSt7collateIwEC2Ey _ZNSt7collateIwEC2Ey .text$_ZNSt7collateIwEC1Ey _ZNSt7collateIwEC1Ey .text$_ZNSt7collateIwEC2EPiy _Z�      NSt7collateIwEC2EPiy .text$_ZNSt7collateIwEC1EPiy _ZNSt7collateIwEC1EPiy .text$_ZNKSt7collateIwE7compareEPKwS2_S2_S2_ _ZNKSt7collateIwE7compareEPKwS2_S2_S2_ .text$_ZNKSt7collateIwE9transformEPKwS2_ _ZNKSt7collateIwE9transformEPKwS2_ .text$_ZNKSt7collateIwE4hashEPKwS2_ _ZNKSt7collateIwE4hashEPKwS2_ .text$_ZNSt7collateIwED2Ev _ZNSt7collateIwED2Ev .text$_ZNSt14collate_bynameIwEC2EPKcy _ZNSt14collate_bynameIwEC2EPKcy .rdata$_ZTVSt14collate_bynameIwE .text$_ZNSt14collate_bynameIwEC1EPKcy _ZNSt14collate_bynameIwEC1EPKcy .text$_ZNSt14collate_bynameIwEC2ERKSsy _ZNSt14collate_bynameIwEC2ERKSsy .text$_ZNSt14collate_bynameIwEC1ERKSsy _ZNSt14collate_bynameIwEC1ERKSsy .text$_ZNSt14collate_bynameIwED2Ev _ZNSt14collate_bynameIwED2Ev .text$_ZSt9use_facetISt5ctypeIwEERKT_RKSt6locale _ZSt9use_facetISt5ctypeIwEERKT_RKSt6locale .text$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmPKwSB_ _ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmPKwSB_ �      .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZSt9use_facetISt7codecvtIwciEERKT_RKSt6locale _ZSt9use_facetISt7codecvtIwciEERKT_RKSt6locale .text$_ZSt9use_facetISt7collateIwEERKT_RKSt6locale _ZSt9use_facetISt7collateIwEERKT_RKSt6locale .data$_ZNSt7collateIwE2idE .rdata$_ZTISt7collateIwE .text$_ZSt9use_facetISt8numpunctIwEERKT_RKSt6locale _ZSt9use_facetISt8numpunctIwEERKT_RKSt6locale .data$_ZNSt8numpunctIwE2idE .rdata$_ZTISt8numpunctIwE .text$_ZNSt16__numpunct_cacheIwE8_M_cacheERKSt6locale _ZNSt16__numpunct_cacheIwE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt7num_pu�      tIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt10moneypunctIwLb1EEERKT_RKSt6locale _ZSt9use_facetISt10moneypunctIwLb1EEERKT_RKSt6locale .data$_ZNSt10moneypunctIwLb1EE2idE .rdata$_ZTISt10moneypunctIwLb1EE .text$_ZNSt18__moneypunct_cacheIwLb1EE8_M_cacheERKSt6locale _ZNSt18__moneypunct_cacheIwLb1EE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt10moneypunctIwLb0EEERKT_RKSt6locale _ZSt9use_facetISt10moneypunctIwLb0EEERKT_RKSt�      6locale .data$_ZNSt10moneypunctIwLb0EE2idE .rdata$_ZTISt10moneypunctIwLb0EE .text$_ZNSt18__moneypunct_cacheIwLb0EE8_M_cacheERKSt6locale _ZNSt18__moneypunct_cacheIwLb0EE8_M_cacheERKSt6locale .text$_ZSt9use_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt11__timepunctIwEERKT_RKSt6locale _ZSt9use_facetISt11__timepunctIwEERKT_RKSt6locale .data$_ZNSt11__timepunctIwE2idE .rdata$_ZTISt11__timepun�      ctIwE .text$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPK2tmcc _ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPK2tmcc .text$_ZSt9use_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale _ZSt9use_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .data$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .rdata$_ZTISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .text$_ZSt9use_facetISt8messagesIwEERKT_RKSt6locale _ZSt9use_facetISt8messagesIwEERKT_RKSt6locale .data$_ZNSt8messagesIwE2idE .rdata$_ZTISt8messagesIwE .text$_Z�      St9has_facetISt5ctypeIwEEbRKSt6locale _ZSt9has_facetISt5ctypeIwEEbRKSt6locale .text$_ZSt9has_facetISt7codecvtIwciEEbRKSt6locale _ZSt9has_facetISt7codecvtIwciEEbRKSt6locale .text$_ZSt9has_facetISt7collateIwEEbRKSt6locale _ZSt9has_facetISt7collateIwEEbRKSt6locale .text$_ZSt9has_facetISt8numpunctIwEEbRKSt6locale _ZSt9has_facetISt8numpunctIwEEbRKSt6locale .text$_ZSt9has_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_facetISt10moneypunctIwLb0EEEbRKSt6locale _ZSt9has_facetISt10moneypunctIwLb0EEEbRKSt6locale .text$_ZSt9has_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_fac�      etISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_facetISt11__timepunctIwEEbRKSt6locale _ZSt9has_facetISt11__timepunctIwEEbRKSt6locale .text$_ZSt9has_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale _ZSt9has_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .text$_ZSt9has_facetISt8messagesIwEEbRKSt6locale _ZSt9has_facetISt8messagesIwEEbRKSt6locale .text$_ZSt14__add_groupingIwEPT_S1_S0_PKcyPKS0_S5_ _ZSt14__add_groupingIwEPT_S1_S0_PKcyPKS0_S5_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE14_M_group_floatEPKcywPKwPwS9_Ri _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE14_M_group_floatEPKcywPKwPwS9_Ri .text$_ZNK�      St7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE12_M_group_intEPKcywRSt8ios_basePwS9_Ri _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE12_M_group_intEPKcywRSt8ios_basePwS9_Ri .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewe _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewe .text$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewRKSbIwS2_SaIwEE _ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11cha�      r_traitsIwEEE6do_putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .text$_ZNSt5__padIwSt11char_traitsIwEE6_S_padERSt8ios_basewPwPKwxx _ZNSt5__padIwSt11char_traitsIwEE6_S_padERSt8ios_basewPwPKwxx .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6_M_padEwxRSt8ios_basePwPKwRi _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6_M_padEwxRSt8ios_basePwPKwRi .text$_ZSt13__int_to_charIwmEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZSt13__int_to_charIwmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .text$_ZSt13__int_to_charIwyEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZSt13__int_to_charIwyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .text$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb1EEEclERKSt6locale _ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb1EEEclERKSt6locale .text$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb0EEEclERKSt6locale _ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb0EEEclERKSt6locale .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIlEES3_S3_RSt8ios_basewT_ _ZNKSt7num_putIwSt19ostreambuf_iterato�      rIwSt11char_traitsIwEEE13_M_insert_intIlEES3_S3_RSt8ios_basewT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewl _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewl .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewl _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewl .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewb _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewb .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intImEES3_S3_RSt8ios_basewT_ _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intImEES3_S3_RSt8ios_basewT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewm _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewm .text$_ZNKSt7num_putIwSt19os�      treambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewm _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewm .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIxEES3_S3_RSt8ios_basewT_ _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIxEES3_S3_RSt8ios_basewT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewx _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewx .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewx _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewx .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIyEES3_S3_RSt8ios_basewT_ _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIyEES3_S3_RSt8ios_basewT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewy _ZN�      KSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewy .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPKv _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPKv .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewy _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewy .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIdEES3_S3_RSt8ios_basewcT_ _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIdEES3_S3_RSt8ios_basewcT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewd _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewd .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIeEES3_S3_RSt8ios_basewcT_ _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_i�      nsert_floatIeEES3_S3_RSt8ios_basewcT_ .text$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewe _ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewe .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istre�      ambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKw _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKw .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_tra�      itsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11�      char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwS�      t11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambu�      f_iteratorIwSt11char_traitsIwEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .text$_ZNKSt7num�      _getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZN�      KSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .text$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_I�      os_IostateRSs .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .text$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE _ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE .text$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSC_ _ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSC_ _GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2E�      RKSsy .data$_ZGVNSt10moneypunctIwLb0EE2idE .data$_ZGVNSt10moneypunctIwLb1EE2idE .data$_ZGVNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt8numpunctIwE2idE .data$_ZGVNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt11__timepunctIwE2idE .data$_ZGVNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .data$_ZGVNSt8messagesIwE2idE .data$_ZGVNSt7collateIwE2idE .rdata$_ZTSSt7collateIwE .rdata$_ZTSSt14collate_bynameIwE .rdata$_ZTISt14collate_bynameIwE .rdata$_ZTSSt8numpunctIwE .rdata$_ZTSSt15numpunct_bynameIwE .rdata$_ZTISt15numpunct_bynameIwE .rdata$_ZTSSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt17__timepunct_cacheIwE .rdata$_ZT�      ISt17__timepunct_cacheIwE .rdata$_ZTSSt11__timepunctIwE .rdata$_ZTSSt10moneypunctIwLb1EE .rdata$_ZTSSt10moneypunctIwLb0EE .rdata$_ZTSSt8messagesIwE .rdata$_ZTSSt14codecvt_bynameIwciE .rdata$_ZTISt14codecvt_bynameIwciE .rdata$_ZTSSt17moneypunct_bynameIwLb0EE .rdata$_ZTISt17moneypunct_bynameIwLb0EE .rdata$_ZTSSt17moneypunct_bynameIwLb1EE .rdata$_ZTISt17moneypunct_bynameIwLb1EE .rdata$_ZTSSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTISt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTISt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .rdata$_ZTSSt15messages_bynameIwE .rdata$_ZT�      ISt15messages_bynameIwE .rdata$_ZTVSt21__ctype_abstract_baseIwE .rdata$_ZTVSt23__codecvt_abstract_baseIwciE .rdata$_ZNSt17moneypunct_bynameIwLb1EE4intlE .rdata$_ZNSt17moneypunct_bynameIwLb0EE4intlE .rdata$_ZNSt10moneypunctIwLb1EE4intlE .rdata$_ZNSt10moneypunctIwLb0EE4intlE .xdata$_ZNKSt10moneypunctIwLb0EE16do_decimal_pointEv .pdata$_ZNKSt10moneypunctIwLb0EE16do_decimal_pointEv .xdata$_ZNKSt10moneypunctIwLb0EE16do_thousands_sepEv .pdata$_ZNKSt10moneypunctIwLb0EE16do_thousands_sepEv .xdata$_ZNKSt10moneypunctIwLb0EE14do_frac_digitsEv .pdata$_ZNKSt10moneypunctIwLb0EE14do_frac_digitsEv .xdata$_ZNKSt10moneypunctIwLb0EE13do_pos_formatEv .pdata$_ZNKSt10moneypunctIwLb0EE13do_pos_formatEv .xdata$_ZNKSt10moneypunctIwLb0EE13do_neg_formatEv .pdata$_ZNKSt10moneypunctIwLb0EE13do_neg_formatEv .xdata$_ZNKSt10moneypunctIwLb1EE16do_decimal_pointEv .pdata$_ZNKSt10moneypunctIwLb1EE16do_decimal_pointEv .xdata$_ZNKSt10moneypunctIwLb1EE16do_thousands_sepEv .pdata$_ZNKSt10moneypunctIwLb1EE16do_thousands_sepEv .xdata$_ZNKSt10m�      oneypunctIwLb1EE14do_frac_digitsEv .pdata$_ZNKSt10moneypunctIwLb1EE14do_frac_digitsEv .xdata$_ZNKSt10moneypunctIwLb1EE13do_pos_formatEv .pdata$_ZNKSt10moneypunctIwLb1EE13do_pos_formatEv .xdata$_ZNKSt10moneypunctIwLb1EE13do_neg_formatEv .pdata$_ZNKSt10moneypunctIwLb1EE13do_neg_formatEv .xdata$_ZNSt17moneypunct_bynameIwLb0EED1Ev .pdata$_ZNSt17moneypunct_bynameIwLb0EED1Ev .xdata$_ZNSt17moneypunct_bynameIwLb1EED1Ev .pdata$_ZNSt17moneypunct_bynameIwLb1EED1Ev .xdata$_ZNKSt8numpunctIwE16do_decimal_pointEv .pdata$_ZNKSt8numpunctIwE16do_decimal_pointEv .xdata$_ZNKSt8numpunctIwE16do_thousands_sepEv .pdata$_ZNKSt8numpunctIwE16do_thousands_sepEv .xdata$_ZNSt15numpunct_bynameIwED1Ev .pdata$_ZNSt15numpunct_bynameIwED1Ev .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13do_date_orderEv .xdata$_ZNKSt8messagesIwE7do_openERKSsRKSt6locale .pdata$_ZNKSt8messagesIwE7do_openERKSsRKSt6locale .xdata$_ZNKSt8messagesIwE8�      do_closeEi .pdata$_ZNKSt8messagesIwE8do_closeEi .xdata$_ZNKSt7collateIwE7do_hashEPKwS2_ .pdata$_ZNKSt7collateIwE7do_hashEPKwS2_ .xdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt17__timepunct_cacheIwED1Ev .pdata$_ZNSt17__timepunct_cacheIwED1Ev .xdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$�      _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED1Ev .xdata$_ZNSt17moneypunct_bynameIwLb0EED0Ev .pdata$_ZNSt17moneypunct_bynameIwLb0EED0Ev .xdata$_ZNSt17moneypunct_bynameIwLb1EED0Ev .pdata$_ZNSt17moneypunct_bynameIwLb1EED0Ev .xdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt15numpunct_bynameIwED0Ev .pdata$_ZNSt15numpunct_bynameIwED0Ev .xdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt�      7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt17__timepunct_cacheIwED0Ev .pdata$_ZNSt17__timepunct_cacheIwED0Ev .xdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED0Ev .xdata$_ZNKSt10moneypunctIwLb0EE11do_groupingEv .pdata$_ZNKSt10moneypunctIwLb0EE11do_groupingEv .xdata$_ZNKSt10moneypu�      nctIwLb1EE11do_groupingEv .pdata$_ZNKSt10moneypunctIwLb1EE11do_groupingEv .xdata$_ZNKSt8numpunctIwE11do_groupingEv .pdata$_ZNKSt8numpunctIwE11do_groupingEv .xdata$_ZNKSt10moneypunctIwLb0EE14do_curr_symbolEv .pdata$_ZNKSt10moneypunctIwLb0EE14do_curr_symbolEv .xdata$_ZNKSt10moneypunctIwLb0EE16do_positive_signEv .pdata$_ZNKSt10moneypunctIwLb0EE16do_positive_signEv .xdata$_ZNKSt10moneypunctIwLb0EE16do_negative_signEv .pdata$_ZNKSt10moneypunctIwLb0EE16do_negative_signEv .xdata$_ZNKSt10moneypunctIwLb1EE14do_curr_symbolEv .pdata$_ZNKSt10moneypunctIwLb1EE14do_curr_symbolEv .xdata$_ZNKSt10moneypunctIwLb1EE16do_positive_signEv .pdata$_ZNKSt10moneypunctIwLb1EE16do_positive_signEv .xdata$_ZNKSt10moneypunctIwLb1EE16do_negative_signEv .pdata$_ZNKSt10moneypunctIwLb1EE16do_negative_signEv .xdata$_ZNKSt8numpunctIwE11do_truenameEv .pdata$_ZNKSt8numpunctIwE11do_truenameEv .xdata$_ZNKSt8numpunctIwE12do_falsenameEv .pdata$_ZNKSt8numpunctIwE12do_falsenameEv .xdata$_ZNSt8messagesIwED1Ev .pdata$_ZNSt8messagesIwED1Ev .xdata$_�      ZNSt8messagesIwED0Ev .pdata$_ZNSt8messagesIwED0Ev .xdata$_ZNSt7collateIwED1Ev .pdata$_ZNSt7collateIwED1Ev .xdata$_ZNSt7collateIwED0Ev .pdata$_ZNSt7collateIwED0Ev .xdata$_ZNSt15messages_bynameIwED1Ev .pdata$_ZNSt15messages_bynameIwED1Ev .xdata$_ZNSt15messages_bynameIwED0Ev .pdata$_ZNSt15messages_bynameIwED0Ev .xdata$_ZNSt14collate_bynameIwED1Ev .pdata$_ZNSt14collate_bynameIwED1Ev .xdata$_ZNSt14collate_bynameIwED0Ev .pdata$_ZNSt14collate_bynameIwED0Ev .xdata$_ZNSt11__timepunctIwED1Ev .pdata$_ZNSt11__timepunctIwED1Ev .xdata$_ZNSt11__timepunctIwED0Ev .pdata$_ZNSt11__timepunctIwED0Ev .xdata$_ZNSt14codecvt_bynameIwciED1Ev .pdata$_ZNSt14codecvt_bynameIwciED1Ev .xdata$_ZNSt14codecvt_bynameIwciED0Ev .pdata$_ZNSt14codecvt_bynameIwciED0Ev .text$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.43 .xdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.43 .pdata$_ZNKSt19istreambuf_iteratorIwSt11char_traitsIwEE6_M_getEv.isra.43 .xdata$_ZNKSt7collateIwE12do_transformEPKwS2_ .pdata$_ZNKSt7�      collateIwE12do_transformEPKwS2_ .xdata$_ZNKSt7collateIwE10do_compareEPKwS2_S2_S2_ .pdata$_ZNKSt7collateIwE10do_compareEPKwS2_S2_S2_ .xdata$_ZNSt18__moneypunct_cacheIwLb0EEC2Ey .pdata$_ZNSt18__moneypunct_cacheIwLb0EEC2Ey .xdata$_ZNSt18__moneypunct_cacheIwLb0EEC1Ey .pdata$_ZNSt18__moneypunct_cacheIwLb0EEC1Ey .xdata$_ZNSt18__moneypunct_cacheIwLb0EED2Ev .pdata$_ZNSt18__moneypunct_cacheIwLb0EED2Ev .xdata$_ZNSt18__moneypunct_cacheIwLb1EEC2Ey .pdata$_ZNSt18__moneypunct_cacheIwLb1EEC2Ey .xdata$_ZNSt18__moneypunct_cacheIwLb1EEC1Ey .pdata$_ZNSt18__moneypunct_cacheIwLb1EEC1Ey .xdata$_ZNSt18__moneypunct_cacheIwLb1EED2Ev .pdata$_ZNSt18__moneypunct_cacheIwLb1EED2Ev .xdata$_ZNSt10moneypunctIwLb0EEC2Ey .pdata$_ZNSt10moneypunctIwLb0EEC2Ey .xdata$_ZNSt10moneypunctIwLb0EEC1Ey .pdata$_ZNSt10moneypunctIwLb0EEC1Ey .xdata$_ZNSt10moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .pdata$_ZNSt10moneypunctIwLb0EEC2EPSt18__moneypunct_cacheIwLb0EEy .xdata$_ZNSt10moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy .pdata$_ZNSt10�      moneypunctIwLb0EEC1EPSt18__moneypunct_cacheIwLb0EEy .xdata$_ZNSt10moneypunctIwLb0EEC2EPiPKcy .pdata$_ZNSt10moneypunctIwLb0EEC2EPiPKcy .xdata$_ZNSt10moneypunctIwLb0EEC1EPiPKcy .pdata$_ZNSt10moneypunctIwLb0EEC1EPiPKcy .xdata$_ZNKSt10moneypunctIwLb0EE13decimal_pointEv .pdata$_ZNKSt10moneypunctIwLb0EE13decimal_pointEv .xdata$_ZNKSt10moneypunctIwLb0EE13thousands_sepEv .pdata$_ZNKSt10moneypunctIwLb0EE13thousands_sepEv .xdata$_ZNKSt10moneypunctIwLb0EE8groupingEv .pdata$_ZNKSt10moneypunctIwLb0EE8groupingEv .xdata$_ZNKSt10moneypunctIwLb0EE11curr_symbolEv .pdata$_ZNKSt10moneypunctIwLb0EE11curr_symbolEv .xdata$_ZNKSt10moneypunctIwLb0EE13positive_signEv .pdata$_ZNKSt10moneypunctIwLb0EE13positive_signEv .xdata$_ZNKSt10moneypunctIwLb0EE13negative_signEv .pdata$_ZNKSt10moneypunctIwLb0EE13negative_signEv .xdata$_ZNKSt10moneypunctIwLb0EE11frac_digitsEv .pdata$_ZNKSt10moneypunctIwLb0EE11frac_digitsEv .xdata$_ZNKSt10moneypunctIwLb0EE10pos_formatEv .pdata$_ZNKSt10moneypunctIwLb0EE10pos_formatEv .xdata$_ZNKSt10moneypunctI�      wLb0EE10neg_formatEv .pdata$_ZNKSt10moneypunctIwLb0EE10neg_formatEv .xdata$_ZNSt10moneypunctIwLb1EEC2Ey .pdata$_ZNSt10moneypunctIwLb1EEC2Ey .xdata$_ZNSt10moneypunctIwLb1EEC1Ey .pdata$_ZNSt10moneypunctIwLb1EEC1Ey .xdata$_ZNSt10moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .pdata$_ZNSt10moneypunctIwLb1EEC2EPSt18__moneypunct_cacheIwLb1EEy .xdata$_ZNSt10moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .pdata$_ZNSt10moneypunctIwLb1EEC1EPSt18__moneypunct_cacheIwLb1EEy .xdata$_ZNSt10moneypunctIwLb1EEC2EPiPKcy .pdata$_ZNSt10moneypunctIwLb1EEC2EPiPKcy .xdata$_ZNSt10moneypunctIwLb1EEC1EPiPKcy .pdata$_ZNSt10moneypunctIwLb1EEC1EPiPKcy .xdata$_ZNKSt10moneypunctIwLb1EE13decimal_pointEv .pdata$_ZNKSt10moneypunctIwLb1EE13decimal_pointEv .xdata$_ZNKSt10moneypunctIwLb1EE13thousands_sepEv .pdata$_ZNKSt10moneypunctIwLb1EE13thousands_sepEv .xdata$_ZNKSt10moneypunctIwLb1EE8groupingEv .pdata$_ZNKSt10moneypunctIwLb1EE8groupingEv .xdata$_ZNKSt10moneypunctIwLb1EE11curr_symbolEv .pdata$_ZNKSt10moneypunctIwLb1EE11curr_s�      ymbolEv .xdata$_ZNKSt10moneypunctIwLb1EE13positive_signEv .pdata$_ZNKSt10moneypunctIwLb1EE13positive_signEv .xdata$_ZNKSt10moneypunctIwLb1EE13negative_signEv .pdata$_ZNKSt10moneypunctIwLb1EE13negative_signEv .xdata$_ZNKSt10moneypunctIwLb1EE11frac_digitsEv .pdata$_ZNKSt10moneypunctIwLb1EE11frac_digitsEv .xdata$_ZNKSt10moneypunctIwLb1EE10pos_formatEv .pdata$_ZNKSt10moneypunctIwLb1EE10pos_formatEv .xdata$_ZNKSt10moneypunctIwLb1EE10neg_formatEv .pdata$_ZNKSt10moneypunctIwLb1EE10neg_formatEv .xdata$_ZNSt17moneypunct_bynameIwLb0EEC2EPKcy .pdata$_ZNSt17moneypunct_bynameIwLb0EEC2EPKcy .xdata$_ZNSt17moneypunct_bynameIwLb0EEC1EPKcy .pdata$_ZNSt17moneypunct_bynameIwLb0EEC1EPKcy .xdata$_ZNSt17moneypunct_bynameIwLb0EEC2ERKSsy .pdata$_ZNSt17moneypunct_bynameIwLb0EEC2ERKSsy .xdata$_ZNSt17moneypunct_bynameIwLb0EEC1ERKSsy .pdata$_ZNSt17moneypunct_bynameIwLb0EEC1ERKSsy .xdata$_ZNSt17moneypunct_bynameIwLb0EED2Ev .pdata$_ZNSt17moneypunct_bynameIwLb0EED2Ev .xdata$_ZNSt17moneypunct_bynameIwLb1EEC2EPKcy .pdata$_ZNSt17moneyp�      unct_bynameIwLb1EEC2EPKcy .xdata$_ZNSt17moneypunct_bynameIwLb1EEC1EPKcy .pdata$_ZNSt17moneypunct_bynameIwLb1EEC1EPKcy .xdata$_ZNSt17moneypunct_bynameIwLb1EEC2ERKSsy .pdata$_ZNSt17moneypunct_bynameIwLb1EEC2ERKSsy .xdata$_ZNSt17moneypunct_bynameIwLb1EEC1ERKSsy .pdata$_ZNSt17moneypunct_bynameIwLb1EEC1ERKSsy .xdata$_ZNSt17moneypunct_bynameIwLb1EED2Ev .pdata$_ZNSt17moneypunct_bynameIwLb1EED2Ev .xdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_�      Ios_IostateRSbIwS2_SaIwEE .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE .xdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewe .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewe .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .xdata$_ZNSt9mon�      ey_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt16__numpunct_cacheIwEC2Ey .pdata$_ZNSt16__numpunct_cacheIwEC2Ey .xdata$_ZNSt16__numpunct_cacheIwEC1Ey .pdata$_ZNSt16__numpunct_cacheIwEC1Ey .xdata$_ZNSt16__numpunct_cacheIwED2Ev .pdata$_ZNSt16__numpunct_cacheIwED2Ev .xdata$_ZNSt8numpunctIwEC2Ey .pdata$_ZNSt8numpunctIwEC2Ey .xdata$_ZNSt8numpunctIwEC1Ey .pdata$_ZNSt8numpunctIwEC1Ey .xdata$_ZNSt8numpunctIwEC2EPSt16__numpunct_cacheIwEy .pdata$_ZNSt8numpunctIwEC2EPSt16__numpunct_cacheIwEy .xdata$_ZNSt8numpunctIwEC1EPSt16__numpunct_cacheIwEy .pdata$_ZNSt8numpunctIwEC1EPSt16__numpunct_cacheIwEy .xdata$_ZNSt8numpunctIwEC2EPiy .pdata$_ZNSt8numpunctIwEC2EPiy .xdata$_ZNSt8numpunctIwEC1EPiy .pdata$_ZNSt8numpunctIwEC1EPiy .xdata$_ZNKSt8numpunctIwE13decimal_pointEv .pdata$_ZNKSt8numpunctIwE13decimal_pointEv .xdata$_ZNKSt8numpunctIwE13thousands_sepEv .pdata$_ZNKSt8numpunctIwE13thousands_sepEv .xdata$_ZNKSt8numpunctIwE8groupi�      ngEv .pdata$_ZNKSt8numpunctIwE8groupingEv .xdata$_ZNKSt8numpunctIwE8truenameEv .pdata$_ZNKSt8numpunctIwE8truenameEv .xdata$_ZNKSt8numpunctIwE9falsenameEv .pdata$_ZNKSt8numpunctIwE9falsenameEv .xdata$_ZNSt15numpunct_bynameIwEC2EPKcy .pdata$_ZNSt15numpunct_bynameIwEC2EPKcy .xdata$_ZNSt15numpunct_bynameIwEC1EPKcy .pdata$_ZNSt15numpunct_bynameIwEC1EPKcy .xdata$_ZNSt15numpunct_bynameIwEC2ERKSsy .pdata$_ZNSt15numpunct_bynameIwEC2ERKSsy .xdata$_ZNSt15numpunct_bynameIwEC1ERKSsy .pdata$_ZNSt15numpunct_bynameIwEC1ERKSsy .xdata$_ZNSt15numpunct_bynameIwED2Ev .pdata$_ZNSt15numpunct_bynameIwED2Ev .xdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .pdata$_ZNKSt7num_getIwSt19�      istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .xdata$_ZNSt7num_getIwSt19istreambuf_itera�      torIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewb .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewb .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewd .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewd .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewe .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewe .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8�      ios_basewPKv .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPKv .xdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt11__timepunctIwEC2Ey .pdata$_ZNSt11__timepunctIwEC2Ey .xdata$_ZNSt11__timepunctIwEC1Ey .pdata$_ZNSt11__timepunctIwEC1Ey .xdata$_ZNSt11__timepunctIwEC2EPSt17__timepunct_cacheIwEy .pdata$_ZNSt11__timepunctIwEC2EPSt17__timepunct_cacheIwEy .xdata$_ZNSt11__timepunctIwEC1EPSt17__timepunct_cacheIwEy .pdata$_ZNSt11__timepunctIwEC1EPSt17__timepunct_cacheIwEy .xdata$_ZNSt11__timepunctIwEC2EPiPKcy .pdata$_ZNSt11__timepunctIwEC2EPiPKcy .xdata$_ZNSt11__timepunctIwEC1EPiPKcy .pdata$_ZNSt11__timepunctIwEC1EPiPKcy .xdata$_ZNKSt11__timepunctIwE15_M_date_formatsEPPKw .pdata$_ZNKSt11__timepunctIwE15_M_date_formatsEPPKw .xdata$_ZNKSt11__timepunctIwE15_M_time_formatsEPPKw .pdata$_ZNKSt11__timepunctIwE15_M_time_formatsEPPKw .xdata$_ZNKSt11__timepunctIwE20_M_date_tim�      e_formatsEPPKw .pdata$_ZNKSt11__timepunctIwE20_M_date_time_formatsEPPKw .xdata$_ZNKSt11__timepunctIwE15_M_am_pm_formatEPKw .pdata$_ZNKSt11__timepunctIwE15_M_am_pm_formatEPKw .xdata$_ZNKSt11__timepunctIwE8_M_am_pmEPPKw .pdata$_ZNKSt11__timepunctIwE8_M_am_pmEPPKw .xdata$_ZNKSt11__timepunctIwE7_M_daysEPPKw .pdata$_ZNKSt11__timepunctIwE7_M_daysEPPKw .xdata$_ZNKSt11__timepunctIwE19_M_days_abbreviatedEPPKw .pdata$_ZNKSt11__timepunctIwE19_M_days_abbreviatedEPPKw .xdata$_ZNKSt11__timepunctIwE9_M_monthsEPPKw .pdata$_ZNKSt11__timepunctIwE9_M_monthsEPPKw .xdata$_ZNKSt11__timepunctIwE21_M_months_abbreviatedEPPKw .pdata$_ZNKSt11__timepunctIwE21_M_months_abbreviatedEPPKw .xdata$_ZNSt11__timepunctIwED2Ev .pdata$_ZNSt11__timepunctIwED2Ev .xdata$_ZNSt17__timepunct_cacheIwEC2Ey .pdata$_ZNSt17__timepunct_cacheIwEC2Ey .xdata$_ZNSt17__timepunct_cacheIwEC1Ey .pdata$_ZNSt17__timepunct_cacheIwEC1Ey .xdata$_ZNSt17__timepunct_cacheIwED2Ev .pdata$_ZNSt17__timepunct_cacheIwED2Ev .xdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt�      11char_traitsIwEEEC2Ey .pdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmcc .pdata$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmcc .xdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .pdata$_ZNS�      t15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .xdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .pdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2Ey .xdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .pdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1Ey .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10date_orderEv .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19ist�      reambuf_iteratorIwSt11char_traitsIwEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE8get_y�      earES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2EPKcy .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1EPKcy .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC2ERKSsy .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEC1ERKSsy .xdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEED2Ev .pdata$_ZNSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_trai�      tsIwEEED2Ev .xdata$_ZNSt8messagesIwEC2Ey .pdata$_ZNSt8messagesIwEC2Ey .xdata$_ZNSt8messagesIwEC1Ey .pdata$_ZNSt8messagesIwEC1Ey .xdata$_ZNSt8messagesIwEC2EPiPKcy .pdata$_ZNSt8messagesIwEC2EPiPKcy .xdata$_ZNSt8messagesIwEC1EPiPKcy .pdata$_ZNSt8messagesIwEC1EPiPKcy .xdata$_ZNKSt8messagesIwE4openERKSsRKSt6locale .pdata$_ZNKSt8messagesIwE4openERKSsRKSt6locale .xdata$_ZNKSt8messagesIwE4openERKSsRKSt6localePKc .pdata$_ZNKSt8messagesIwE4openERKSsRKSt6localePKc .xdata$_ZNKSt8messagesIwE3getEiiiRKSbIwSt11char_traitsIwESaIwEE .pdata$_ZNKSt8messagesIwE3getEiiiRKSbIwSt11char_traitsIwESaIwEE .xdata$_ZNKSt8messagesIwE5closeEi .pdata$_ZNKSt8messagesIwE5closeEi .xdata$_ZNSt8messagesIwED2Ev .pdata$_ZNSt8messagesIwED2Ev .xdata$_ZNKSt8messagesIwE18_M_convert_to_charERKSbIwSt11char_traitsIwESaIwEE .pdata$_ZNKSt8messagesIwE18_M_convert_to_charERKSbIwSt11char_traitsIwESaIwEE .xdata$_ZNKSt8messagesIwE20_M_convert_from_charEPc .pdata$_ZNKSt8messagesIwE20_M_convert_from_charEPc .xdata$_ZNSt15messages_bynameIwEC2EPKcy .pdata$_�      ZNSt15messages_bynameIwEC2EPKcy .xdata$_ZNSt15messages_bynameIwEC1EPKcy .pdata$_ZNSt15messages_bynameIwEC1EPKcy .xdata$_ZNSt15messages_bynameIwEC2ERKSsy .pdata$_ZNSt15messages_bynameIwEC2ERKSsy .xdata$_ZNSt15messages_bynameIwEC1ERKSsy .pdata$_ZNSt15messages_bynameIwEC1ERKSsy .xdata$_ZNSt15messages_bynameIwED2Ev .pdata$_ZNSt15messages_bynameIwED2Ev .text$_ZNSt12ctype_bynameIwEC2ERKSsy .xdata$_ZNSt12ctype_bynameIwEC2ERKSsy .pdata$_ZNSt12ctype_bynameIwEC2ERKSsy .xdata$_ZNSt14codecvt_bynameIwciEC2EPKcy .pdata$_ZNSt14codecvt_bynameIwciEC2EPKcy .xdata$_ZNSt14codecvt_bynameIwciEC1EPKcy .pdata$_ZNSt14codecvt_bynameIwciEC1EPKcy .xdata$_ZNSt14codecvt_bynameIwciEC2ERKSsy .pdata$_ZNSt14codecvt_bynameIwciEC2ERKSsy .xdata$_ZNSt14codecvt_bynameIwciEC1ERKSsy .pdata$_ZNSt14codecvt_bynameIwciEC1ERKSsy .xdata$_ZNSt14codecvt_bynameIwciED2Ev .pdata$_ZNSt14codecvt_bynameIwciED2Ev .xdata$_ZNSt7collateIwEC2Ey .pdata$_ZNSt7collateIwEC2Ey .xdata$_ZNSt7collateIwEC1Ey .pdata$_ZNSt7collateIwEC1Ey .xdata$_ZNSt7collateIwEC2EPiy .pd�      ata$_ZNSt7collateIwEC2EPiy .xdata$_ZNSt7collateIwEC1EPiy .pdata$_ZNSt7collateIwEC1EPiy .xdata$_ZNKSt7collateIwE7compareEPKwS2_S2_S2_ .pdata$_ZNKSt7collateIwE7compareEPKwS2_S2_S2_ .xdata$_ZNKSt7collateIwE9transformEPKwS2_ .pdata$_ZNKSt7collateIwE9transformEPKwS2_ .xdata$_ZNKSt7collateIwE4hashEPKwS2_ .pdata$_ZNKSt7collateIwE4hashEPKwS2_ .xdata$_ZNSt7collateIwED2Ev .pdata$_ZNSt7collateIwED2Ev .xdata$_ZNSt14collate_bynameIwEC2EPKcy .pdata$_ZNSt14collate_bynameIwEC2EPKcy .xdata$_ZNSt14collate_bynameIwEC1EPKcy .pdata$_ZNSt14collate_bynameIwEC1EPKcy .xdata$_ZNSt14collate_bynameIwEC2ERKSsy .pdata$_ZNSt14collate_bynameIwEC2ERKSsy .xdata$_ZNSt14collate_bynameIwEC1ERKSsy .pdata$_ZNSt14collate_bynameIwEC1ERKSsy .xdata$_ZNSt14collate_bynameIwED2Ev .pdata$_ZNSt14collate_bynameIwED2Ev .xdata$_ZSt9use_facetISt5ctypeIwEERKT_RKSt6locale .pdata$_ZSt9use_facetISt5ctypeIwEERKT_RKSt6locale .xdata$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmPKwSB_ .pdata$_ZNKSt8time_putIwSt19ostre�      ambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewPK2tmPKwSB_ .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_numES3_S3_RiiiyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZSt9use_facetISt7codecvtIwciEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7codecvtIwciEERKT_RKSt6locale .xdata$_ZSt9use_facetISt7collateIwEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7collateIwEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8numpunctIwEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8numpunctIwEERKT_RKSt6locale .xdata$_ZNSt16__numpunct_cacheIwE8_M_cacheERKSt6locale .pdata$_ZNSt16__numpunct_cacheIwE8_M_cacheERKSt6locale .xdata$_ZSt9use_fac�      etISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt10moneypunctIwLb1EEERKT_RKSt6locale .pdata$_ZSt9use_facetISt10moneypunctIwLb1EEERKT_RKSt6locale .xdata$_ZNSt18__moneypunct_cacheIwLb1EE8_M_cacheERKSt6locale .pdata$_ZNSt18__moneypunct_cacheIwLb1EE8_M_cacheERKSt6locale .xdata$_ZSt9use_facetISt10moneypunctIwLb0EEERKT_RKSt6locale .pdata$_ZSt9use_facetISt10moneypunctIwLb0EEERKT_RKSt6locale .xdata$_ZNSt18__moneypunct_cacheIwLb0EE8_M_cacheERKSt6locale .pdata$_ZNSt18__moneypunct_cacheIwLb0EE8_M_cacheERKSt6locale .xdata$_ZSt9use_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char�      _traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt11__timepunctIwEERKT_RKSt6locale .pdata$_ZSt9use_facetISt11__timepunctIwEERKT_RKSt6locale .xdata$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPK2tmcc .pdata$_ZNKSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPK2tmcc .xdata$_ZSt9use_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEERKT_RKSt6locale .xdata$_ZSt9use_facetISt8messagesIwEERKT_RKSt6locale .pdata$_ZSt9use_facetISt8messagesI�      wEERKT_RKSt6locale .xdata$_ZSt9has_facetISt5ctypeIwEEbRKSt6locale .pdata$_ZSt9has_facetISt5ctypeIwEEbRKSt6locale .xdata$_ZSt9has_facetISt7codecvtIwciEEbRKSt6locale .pdata$_ZSt9has_facetISt7codecvtIwciEEbRKSt6locale .xdata$_ZSt9has_facetISt7collateIwEEbRKSt6locale .pdata$_ZSt9has_facetISt7collateIwEEbRKSt6locale .xdata$_ZSt9has_facetISt8numpunctIwEEbRKSt6locale .pdata$_ZSt9has_facetISt8numpunctIwEEbRKSt6locale .xdata$_ZSt9has_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt10moneypunctIwLb0EEEbRKSt6locale .pdata$_ZSt9has_facetISt10moneypunctIwLb0EEEbRKSt6locale .xdata$_ZSt9has_facetISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetI�      St9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt11__timepunctIwEEbRKSt6locale .pdata$_ZSt9has_facetISt11__timepunctIwEEbRKSt6locale .xdata$_ZSt9has_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .pdata$_ZSt9has_facetISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEEbRKSt6locale .xdata$_ZSt9has_facetISt8messagesIwEEbRKSt6locale .pdata$_ZSt9has_facetISt8messagesIwEEbRKSt6locale .xdata$_ZSt14__add_groupingIwEPT_S1_S0_PKcyPKS0_S5_ .pdata$_ZSt14__add_groupingIwEPT_S1_S0_PKcyPKS0_S5_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIw�      EEE14_M_group_floatEPKcywPKwPwS9_Ri .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE14_M_group_floatEPKcywPKwPwS9_Ri .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE12_M_group_intEPKcywRSt8ios_basePwS9_Ri .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE12_M_group_intEPKcywRSt8ios_basePwS9_Ri .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb1EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE9_M_insertILb0EEES3_S3_RSt8ios_basewRKSbIwS2_SaIwEE .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewe .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putE�      S3_bRSt8ios_basewe .xdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .pdata$_ZNKSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_bRSt8ios_basewRKSbIwS2_SaIwEE .xdata$_ZNSt5__padIwSt11char_traitsIwEE6_S_padERSt8ios_basewPwPKwxx .pdata$_ZNSt5__padIwSt11char_traitsIwEE6_S_padERSt8ios_basewPwPKwxx .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6_M_padEwxRSt8ios_basePwPKwRi .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6_M_padEwxRSt8ios_basePwPKwRi .xdata$_ZSt13__int_to_charIwmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .pdata$_ZSt13__int_to_charIwmEiPT_T0_PKS0_St13_Ios_Fmtflagsb .xdata$_ZSt13__int_to_charIwyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .pdata$_ZSt13__int_to_charIwyEiPT_T0_PKS0_St13_Ios_Fmtflagsb .xdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb1EEEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb1EEEclERKSt6locale .xdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb0E�      EEclERKSt6locale .pdata$_ZNKSt11__use_cacheISt18__moneypunct_cacheIwLb0EEEclERKSt6locale .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIlEES3_S3_RSt8ios_basewT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIlEES3_S3_RSt8ios_basewT_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewl .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewl .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewl .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewl .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewb .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewb .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intImEES3_S3_RSt8ios_basewT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iter�      atorIwSt11char_traitsIwEEE13_M_insert_intImEES3_S3_RSt8ios_basewT_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewm .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewm .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewm .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewm .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIxEES3_S3_RSt8ios_basewT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIxEES3_S3_RSt8ios_basewT_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewx .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewx .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewx .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8io�      s_basewx .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIyEES3_S3_RSt8ios_basewT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE13_M_insert_intIyEES3_S3_RSt8ios_basewT_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewy .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewy .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPKv .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewPKv .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewy .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE3putES3_RSt8ios_basewy .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIdEES3_S3_RSt8ios_basewcT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIdEES3_S3_RSt8ios_basewcT_ .xd�      ata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewd .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewd .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIeEES3_S3_RSt8ios_basewcT_ .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE15_M_insert_floatIeEES3_S3_RSt8ios_basewcT_ .xdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewe .pdata$_ZNKSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE6do_putES3_RSt8ios_basewe .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE15_M_extract_nameES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .pdata$_ZNKSt8time_g�      etIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE24_M_extract_wday_or_monthES3_S3_RiPPKwyRSt8ios_baseRSt12_Ios_Iostate .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKw .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKw .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_Iostat�      eP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmcc .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt7num_getIwSt19istreambuf_iterato�      rIwSt11char_traitsIwEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_Io�      stateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6�      do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .pdata$_ZNKSt7num_getIwSt19istreambu�      f_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIxEES3_S3_S3_RSt8�      ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwS�      t11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv .xdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .pdata$_ZNKSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8�      ios_baseRSt12_Ios_IostateRe .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe .xdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE .pdata$_ZNKSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSbIwS2_SaIwEE .xdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSC_ .pdata$_ZNKSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKwSC_ .text.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKSsy .xdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKSsy .pdata.startup._GLOBAL__sub_I__ZNSt12ctype_bynameIwEC2ERKSsy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEPw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEPw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESa�      IwEE9_M_lengthEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_lengthEy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_capacityEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_capacityEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_set_lengthEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_set_lengthEy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_is_localEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_is_localEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_�      M_createERyy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_createERyy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_disposeEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_disposeEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_destroyEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_destroyEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE18_M_construct_aux_2Eyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE18_M_construct_aux_2Eyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .text$_ZNKSt7__cxx1112basic_strin 	      gIwSt11char_traitsIwESaIwEE8_M_checkEyPKc _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_limitEyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_limitEyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_copyEPwPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_copyEPwPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_moveEPwPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_moveEPwPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_S_assignEPwyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_S_assignEPwyw .text$_ZNSt7__cxx1112	      basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS4_EESA_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS4_EESA_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS5_S5_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS5_S5_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS7_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS7_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_S_compareEyy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_S_compareEyy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_assignERKS4_ _ZNSt7__cxx1112basic_stri	      ngIwSt11char_traitsIwESaIwEE9_M_assignERKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_mutateEyyPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_mutateEyyPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_eraseEyy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_eraseEyy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2Ev _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2Ev .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1Ev _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1Ev .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EywRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EywRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_tra	      itsIwESaIwEEC1EywRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EywRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED2Ev _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED2Ev .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED1Ev _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED1Ev .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSERKS4_ .text$_ZNSt7__cxx1112ba	      sic_stringIwSt11char_traitsIwESaIwEEaSEOS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEOS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .	      text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6cbeginEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6cbeginEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4cendEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4cendEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7crbeginEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7crbeginEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5crendEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5crendEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4sizeEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4sizeEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6lengthEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6lengthEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8max_sizeEv _ZNKSt7__cxx1112bas	      ic_stringIwSt11char_traitsIwESaIwEE8max_sizeEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8capacityEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8capacityEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7reserveEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7reserveEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13shrink_to_fitEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5clearEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5clearEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5emptyEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5emptyEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .text$_ZNKSt7__cxx1112basic_stringIwSt11c	      har_traitsIwESaIwEE2atEy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9push_backEw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9push_backEw .text$_ZNSt7__cxx1112basic_	      stringIwSt11char_traitsIwESaIwEE6assignERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEOS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEOS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEyy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEyy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8pop_backEv _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8pop_backEv .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyy		      w _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEw _ZNSt7__cxx1112basic_stringIwSt11char_t
	      raitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_yw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_yw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_replaceEyyPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_replaceEyyPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_yy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKwy _ZNSt7__cxx11	      12basic_stringIwSt11char_traitsIwESaIwEE6assignEPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKwy 	      _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_RKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_RKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_y _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_y .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_yy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_yy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIw	      EE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_PwSA_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_PwSA_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_S8_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_S8_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_St16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_St16initializer_listIwE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EESt16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EESt16initializer_listIwE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_	      EES9_NS6_IPwS4_EESB_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_NS6_IPwS4_EESB_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S9_S9_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S9_S9_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_appendEPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_appendEPKwy .	      text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLERKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_yy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEPKw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEPKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .text$_ZNSt7__cxx1112basic_stringIwSt	      11char_traitsIwESaIwEE6appendESt16initializer_listIwE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4copyEPwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4copyEPwyy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4swapERS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4swapERS4_ .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5c_strEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5c_strEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4dataEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4dataEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13get_allocatorEv _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13get_allocatorEv .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaI	      wEE4findERKS4_y _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindERKS4_y _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofERKS4_y _ZNKSt7__cxx1112basic_string	      IwSt11char_traitsIwESaIwEE13find_first_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofERKS4_y _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .text$_ZNKSt7__cxx1112basic_strin	      gIwSt11char_traitsIwESaIwEE12find_last_ofEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS4_y _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_o	      fERKS4_y _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS4_y .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareERKS4_ _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareERKS4_ .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_ _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_ .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_yy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_yy .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEPKw _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEPKw .text$_ZNKSt7__cxx1112b	      asic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKw _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKw .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKwy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwOS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwOS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwOS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwOS3_ .text$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ _ZStplIwSt11char_tra	      itsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .text$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ _ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvT_SA_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvT_SA_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_const	      ructIN9__gnu_cxx17__normal_iteratorIPKwS4_EEEEvT_SB_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKwS4_EEEEvT_SB_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPwEEvT_S7_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPwEEvT_S7_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_ .text$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx	      1112basic_stringIT_T0_T1_EERKS8_SA_ _ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPwvEET_S7_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPwvEET_S7_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPwvEET_S7_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPwvEET_S7_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPKwEEvT_S8_St20forward_iterator_tag _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPKwEEvT_S8_St20forward_iterator_tag .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yy _ZNSt7__cxx1112basic_stringIwSt11ch	      ar_traitsIwESaIwEEC2ERKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yyRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yyRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yyRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yyRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwyRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwyRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwyRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwyRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwRKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwRKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwRKS3_ .text$_ZNSt7__cxx	      1112basic_stringIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPKwvEET_S8_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPKwvEET_S8_RKS3_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPKwvEET_S8_RKS3_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPKwvEET_S8_RKS3_ .text$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6substrEyy _ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6substrEyy .text$_ZN9__gnu_cxxeqIPwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ _ZN9__gnu_cxxeqIPwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ .text$_ZN9__gnu_c	      xxeqIPKwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ _ZN9__gnu_cxxeqIPKwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ .rdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4nposE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEPw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEPw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_lengthEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_lengthEy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_M_dataEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local_dataEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_local	      _dataEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_capacityEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_capacityEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_set_lengthEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_M_set_lengthEy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_is_localEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_is_localEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_createERyy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_createERyy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_disposeEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_disposeEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_destroyEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_destroyEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructEyw .pdata$_ZNSt7__cxx	      1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE18_M_construct_aux_2Eyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE18_M_construct_aux_2Eyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16_M_get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_checkEyPKc .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE15_M_check_lengthEyyPKc .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_limitEyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_l	      imitEyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE11_M_disjunctEPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_copyEPwPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_copyEPwPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_moveEPwPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7_S_moveEPwPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_S_assignEPwyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_S_assignEPwyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIS5_S4_EES8_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS4_EESA_ .pdata$_ZNSt7__cxx1112basic_str	      ingIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwN9__gnu_cxx17__normal_iteratorIPKwS4_EESA_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS5_S5_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwS5_S5_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS7_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13_S_copy_charsEPwPKwS7_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_S_compareEyy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_S_compareEyy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_assignERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_assignERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_mutateEyyPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_mutateEyyPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8_M_eraseEyy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traits 	      IwESaIwEE8_M_eraseEyy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2Ev .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2Ev .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1Ev .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1Ev .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EywRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EywRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EywRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EywRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt!	      11char_traitsIwESaIwEEC1EOS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EOS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EOS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED2Ev .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED2Ev .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED1Ev .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEED1Ev .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEOS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEOS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv .pdata$_ZNSt7__cxx1112b"	      asic_stringIwSt11char_traitsIwESaIwEE5beginEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5beginEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE3endEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6rbeginEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4rendEv .xda#	      ta$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6cbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6cbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4cendEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4cendEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7crbeginEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7crbeginEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5crendEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5crendEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4sizeEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4sizeEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6lengthEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6lengthEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8max_sizeEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8max_sizeEv .xdata$_ZNKSt7__cxx1112basic_s$	      tringIwSt11char_traitsIwESaIwEE8capacityEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8capacityEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7reserveEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7reserveEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13shrink_to_fitEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5clearEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5clearEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5emptyEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5emptyEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEixEy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2%	      atEy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE2atEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5frontEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4backEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9push_backEw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaI&	      wEE9push_backEw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEOS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEOS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEyy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEyy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE8pop_backEv .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE'	      8pop_backEv .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE14_M_replace_auxEyyyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6resizeEy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyyw (	      .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_yw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_yw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPKwS4_EEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_replaceEyyPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE10_M_replaceEyyPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11ch)	      ar_traitsIwESaIwEE6assignERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSESt16initializer_listIwE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignESt16initializer_listIwE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6assignEPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEaSEPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt1*	      1char_traitsIwESaIwEEaSEPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_RKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_RKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_y .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_y .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEy+	      yRKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyRKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyRKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_PwSA_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_PwSA_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_S8_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_S8_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_St16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_St16initializer_listIwE .xdata$_ZNSt7__cxx1112basic_string,	      IwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EESt16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EESt16initializer_listIwE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_NS6_IPwS4_EESB_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_NS6_IPwS4_EESB_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S9_S9_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S9_S9_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEyPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEyyPKw .xda-	      ta$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPKwS4_EES9_S8_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_appendEPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE9_M_appendEPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwE.	      SaIwEE6appendEPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendEPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEPKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLEPKw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEpLESt16initializer_listIwE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6appendESt16initializer_listIwE .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4copyEPwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4copyEPwyy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4swapERS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4swapERS4_ .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5c_strEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5c_strEv .xdata$_/	      ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4dataEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4dataEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13get_allocatorEv .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13get_allocatorEv .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4findEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwyy .x0	      data$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5rfindEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEwy .p1	      data$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE13find_first_ofEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12find_last_ofEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .pdata$_ZNKSt7__cxx1112ba2	      sic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE17find_first_not_ofEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwyy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS4_y .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofERKS4_y .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEPKwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .pdata$_ZNKSt7_3	      _cxx1112basic_stringIwSt11char_traitsIwESaIwEE16find_last_not_ofEwy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareERKS4_ .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareERKS4_ .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_ .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_ .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_yy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyRKS4_yy .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEPKw .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEPKw .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKw .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKw .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKwy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7compareEyyPKwy .xdata$_ZNSt7__cxx1112basi4	      c_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwOS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC2EPwOS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwOS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_Alloc_hiderC1EPwOS3_ .xdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .pdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EEPKS5_RKS8_ .xdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ .pdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EES5_RKS8_ .xdata$_ZNSt7__cxx1112basi5	      c_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvT_SA_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvT_SA_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IN9__gnu_cxx17__normal_iteratorIPwS4_EEvEET_SA_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKwS4_EEEEvT_SB_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIN9__gnu_cxx17__normal_iteratorIPKwS4_EEEEvT_SB_St20forward_iterator_6	      tag .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPwEEvT_S7_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPwEEvT_S7_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_ .xdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .pdata$_ZStplIwSt11char_traitsIwESaIwEENSt7__cxx1112basic_stringIT_T0_T1_EERKS8_SA_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsI7	      wESaIwEEC2IPwvEET_S7_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPwvEET_S7_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPwvEET_S7_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPwvEET_S7_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPKwEEvT_S8_St20forward_iterator_tag .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE12_M_constructIPKwEEvT_S8_St20forward_iterator_tag .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yy .pdata$_ZNSt7__cx8	      x1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ERKS4_yyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ERKS4_yyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwyRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwyRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2EPKwRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwRKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1EPKwRKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ESt16initializer9	      _listIwERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2ESt16initializer_listIwERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1ESt16initializer_listIwERKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPKwvEET_S8_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC2IPKwvEET_S8_RKS3_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPKwvEET_S8_RKS3_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEC1IPKwvEET_S8_RKS3_ .xdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6substrEyy .pdata$_ZNKSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6substrEyy .xdata$_ZN9__gnu_cxxeqIPwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ .pdata$_ZN9__gnu_cxxeqIPwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESD_ .xdata$_ZN9__gnu_cxxeqIPKwNSt7:	      __cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ .pdata$_ZN9__gnu_cxxeqIPKwNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEEEEEbRKNS_17__normal_iteratorIT_T0_EESE_ _ZNKSt9bad_alloc4whatEv _ZNSt9bad_allocD2Ev .rdata$_ZTVSt9bad_alloc _ZNSt9bad_allocD1Ev _ZNSt9bad_allocD0Ev .text$_ZNKSt9bad_alloc4whatEv .xdata$_ZNKSt9bad_alloc4whatEv .pdata$_ZNKSt9bad_alloc4whatEv .text$_ZNSt9bad_allocD2Ev .xdata$_ZNSt9bad_allocD2Ev .pdata$_ZNSt9bad_allocD2Ev .text$_ZNSt9bad_allocD0Ev .xdata$_ZNSt9bad_allocD0Ev .pdata$_ZNSt9bad_allocD0Ev _ZNKSt8bad_cast4whatEv _ZNSt8bad_castD2Ev .rdata$_ZTVSt8bad_cast _ZNSt8bad_castD1Ev _ZNSt8bad_castD0Ev .text$_ZNKSt8bad_cast4whatEv .xdata$_ZNKSt8bad_cast4whatEv .pdata$_ZNKSt8bad_cast4whatEv .text$_ZNSt8bad_castD2Ev .xdata$_ZNSt8bad_castD2Ev .pdata$_ZNSt8bad_castD2Ev .text$_ZNSt8bad_castD0Ev .xdata$_ZNSt8bad_castD0Ev .pdata$_ZNSt8bad_castD0Ev _ZNKSt10bad_typeid4whatEv _ZNSt10bad_typeidD2Ev .rdata$_ZTVSt10bad_typeid _ZNSt10bad_typeidD1Ev _ZNSt10bad;	      _typeidD0Ev .text$_ZNKSt10bad_typeid4whatEv .xdata$_ZNKSt10bad_typeid4whatEv .pdata$_ZNKSt10bad_typeid4whatEv .text$_ZNSt10bad_typeidD2Ev .xdata$_ZNSt10bad_typeidD2Ev .pdata$_ZNSt10bad_typeidD2Ev .text$_ZNSt10bad_typeidD0Ev .xdata$_ZNSt10bad_typeidD0Ev .pdata$_ZNSt10bad_typeidD0Ev _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PPv _ZNK10__cxxabiv117__class_type_info20__do_find_public_srcExPKvPKS0_S2_ _ZN10__cxxabiv117__class_type_infoD2Ev .rdata$_ZTVN10__cxxabiv117__class_type_infoE _ZN10__cxxabiv117__class_type_infoD1Ev _ZN10__cxxabiv117__class_type_infoD0Ev _ZNK10__cxxabiv117__class_type_info12__do_dyncastExNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE _ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj .rdata$_ZTSSt9type_info .rdata$_ZTISt9type_info .rdata$_ZTSN10__cxxabiv117__class_type_infoE .rdata$_ZTIN10__cxxabiv117__class_type_infoE .text$_ZNK10__cxxabiv117__class_type_info11__do_up<	      castEPKS0_PPv .xdata$_ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PPv .pdata$_ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PPv .text$_ZNK10__cxxabiv117__class_type_info20__do_find_public_srcExPKvPKS0_S2_ .xdata$_ZNK10__cxxabiv117__class_type_info20__do_find_public_srcExPKvPKS0_S2_ .pdata$_ZNK10__cxxabiv117__class_type_info20__do_find_public_srcExPKvPKS0_S2_ .text$_ZN10__cxxabiv117__class_type_infoD2Ev .xdata$_ZN10__cxxabiv117__class_type_infoD2Ev .pdata$_ZN10__cxxabiv117__class_type_infoD2Ev .text$_ZN10__cxxabiv117__class_type_infoD0Ev .xdata$_ZN10__cxxabiv117__class_type_infoD0Ev .pdata$_ZN10__cxxabiv117__class_type_infoD0Ev .text$_ZNK10__cxxabiv117__class_type_info12__do_dyncastExNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE .xdata$_ZNK10__cxxabiv117__class_type_info12__do_dyncastExNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE .pdata$_ZNK10__cxxabiv117__class_type_info12__do_dyncastExNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE .text$_ZNK10__cxxabiv117=	      __class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE .xdata$_ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE .pdata$_ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE .text$_ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj .xdata$_ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj .pdata$_ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj .text$_ZdlPv .xdata$_ZdlPv .pdata$_ZdlPv .text$_ZdlPvy .xdata$_ZdlPvy .pdata$_ZdlPvy .text$_ZdaPv .xdata$_ZdaPv .pdata$_ZdaPv __dynamic_cast .text$__dynamic_cast .xdata$__dynamic_cast .pdata$__dynamic_cast _ZN12_GLOBAL__N_114emergency_poolE _ZN12_GLOBAL__N_14pool4freeEPv.constprop.2 _ZN12_GLOBAL__N_14pool8allocateEy.constprop.3 _ZN9__gnu_cxx9__freeresEv __cxa_free_exception __cxa_allocate_dependent_exception __cxa_free_dependent_exception _GLOBAL__sub_I__ZN9__gnu_cxx9__freeresEv __cxa_allocate_exception .text$_ZN12_GLOBAL__N_14pool4freeEPv.constprop.>	      2 .xdata$_ZN12_GLOBAL__N_14pool4freeEPv.constprop.2 .pdata$_ZN12_GLOBAL__N_14pool4freeEPv.constprop.2 .text$_ZN12_GLOBAL__N_14pool8allocateEy.constprop.3 .xdata$_ZN12_GLOBAL__N_14pool8allocateEy.constprop.3 .pdata$_ZN12_GLOBAL__N_14pool8allocateEy.constprop.3 .text$_ZN9__gnu_cxx9__freeresEv .xdata$_ZN9__gnu_cxx9__freeresEv .pdata$_ZN9__gnu_cxx9__freeresEv .text$__cxa_allocate_exception .xdata$__cxa_allocate_exception .pdata$__cxa_allocate_exception .text$__cxa_free_exception .xdata$__cxa_free_exception .pdata$__cxa_free_exception .text$__cxa_allocate_dependent_exception .xdata$__cxa_allocate_dependent_exception .pdata$__cxa_allocate_dependent_exception .text$__cxa_free_dependent_exception .xdata$__cxa_free_dependent_exception .pdata$__cxa_free_dependent_exception .text.startup._GLOBAL__sub_I__ZN9__gnu_cxx9__freeresEv .xdata.startup._GLOBAL__sub_I__ZN9__gnu_cxx9__freeresEv .pdata.startup._GLOBAL__sub_I__ZN9__gnu_cxx9__freeresEv .data$_ZN12_GLOBAL__N_114emergency_poolE __cxa_bad_cast __cxa_bad_typeid __?	      cxa_throw_bad_array_new_length .rdata$.refptr._ZTVSt20bad_array_new_length .rdata$_ZTISt20bad_array_new_length .rdata$_ZTSSt20bad_array_new_length .rdata$.refptr._ZNSt20bad_array_new_lengthD1Ev .text$__cxa_bad_cast .xdata$__cxa_bad_cast .pdata$__cxa_bad_cast .text$__cxa_bad_typeid .xdata$__cxa_bad_typeid .pdata$__cxa_bad_typeid .text$__cxa_throw_bad_array_new_length .xdata$__cxa_throw_bad_array_new_length .pdata$__cxa_throw_bad_array_new_length __cxa_get_exception_ptr __cxa_begin_catch __cxa_end_catch _ZSt18uncaught_exceptionv _ZSt19uncaught_exceptionsv .text$__cxa_get_exception_ptr .xdata$__cxa_get_exception_ptr .pdata$__cxa_get_exception_ptr .text$__cxa_begin_catch .xdata$__cxa_begin_catch .pdata$__cxa_begin_catch .text$__cxa_end_catch .xdata$__cxa_end_catch .pdata$__cxa_end_catch .text$_ZSt18uncaught_exceptionv .xdata$_ZSt18uncaught_exceptionv .pdata$_ZSt18uncaught_exceptionv .text$_ZSt19uncaught_exceptionsv .xdata$_ZSt19uncaught_exceptionsv .pdata$_ZSt19uncaught_exceptionsv _ZNSt9exceptionD2Ev _ZN@	      St9exceptionD1Ev _ZNSt13bad_exceptionD2Ev _ZNSt13bad_exceptionD1Ev _ZNKSt9exception4whatEv _ZGTtNKSt9exception4whatEv _ZNKSt13bad_exception4whatEv _ZGTtNKSt13bad_exception4whatEv _ZNSt9exceptionD0Ev _ZNSt13bad_exceptionD0Ev _ZN10__cxxabiv115__forced_unwindD2Ev _ZN10__cxxabiv115__forced_unwindD1Ev _ZN10__cxxabiv115__forced_unwindD0Ev _ZN10__cxxabiv119__foreign_exceptionD2Ev _ZN10__cxxabiv119__foreign_exceptionD1Ev _ZN10__cxxabiv119__foreign_exceptionD0Ev _ZGTtNKSt9exceptionD1Ev _ZGTtNKSt13bad_exceptionD1Ev .rdata$_ZTSN10__cxxabiv119__foreign_exceptionE .rdata$_ZTIN10__cxxabiv119__foreign_exceptionE .rdata$_ZTVSt9exception .rdata$_ZTVSt13bad_exception .rdata$_ZTVN10__cxxabiv115__forced_unwindE .rdata$_ZTVN10__cxxabiv119__foreign_exceptionE .text$_ZNSt9exceptionD2Ev .xdata$_ZNSt9exceptionD2Ev .pdata$_ZNSt9exceptionD2Ev .text$_ZNSt13bad_exceptionD2Ev .xdata$_ZNSt13bad_exceptionD2Ev .pdata$_ZNSt13bad_exceptionD2Ev .text$_ZNKSt9exception4whatEv .xdata$_ZNKSt9exception4whatEv .pdata$_ZNKSt9exception4whatEv .A	      text$_ZNKSt13bad_exception4whatEv .xdata$_ZNKSt13bad_exception4whatEv .pdata$_ZNKSt13bad_exception4whatEv .text$_ZNSt9exceptionD0Ev .xdata$_ZNSt9exceptionD0Ev .pdata$_ZNSt9exceptionD0Ev .text$_ZNSt13bad_exceptionD0Ev .xdata$_ZNSt13bad_exceptionD0Ev .pdata$_ZNSt13bad_exceptionD0Ev .text$_ZN10__cxxabiv115__forced_unwindD2Ev .xdata$_ZN10__cxxabiv115__forced_unwindD2Ev .pdata$_ZN10__cxxabiv115__forced_unwindD2Ev .text$_ZN10__cxxabiv115__forced_unwindD0Ev .xdata$_ZN10__cxxabiv115__forced_unwindD0Ev .pdata$_ZN10__cxxabiv115__forced_unwindD0Ev .text$_ZN10__cxxabiv119__foreign_exceptionD2Ev .xdata$_ZN10__cxxabiv119__foreign_exceptionD2Ev .pdata$_ZN10__cxxabiv119__foreign_exceptionD2Ev .text$_ZN10__cxxabiv119__foreign_exceptionD0Ev .xdata$_ZN10__cxxabiv119__foreign_exceptionD0Ev .pdata$_ZN10__cxxabiv119__foreign_exceptionD0Ev .text$_ZGTtNKSt9exceptionD1Ev .xdata$_ZGTtNKSt9exceptionD1Ev .pdata$_ZGTtNKSt9exceptionD1Ev .text$_ZGTtNKSt13bad_exceptionD1Ev .xdata$_ZGTtNKSt13bad_exceptionD1Ev .pdata$_ZGTtNKSt13bad_exB	      ceptionD1Ev __cxa_get_globals __emutls_v._ZZN12_GLOBAL__N_110get_globalEvE6global __cxa_get_globals_fast .text$__cxa_get_globals .xdata$__cxa_get_globals .pdata$__cxa_get_globals .text$__cxa_get_globals_fast .xdata$__cxa_get_globals_fast .pdata$__cxa_get_globals_fast .data$__emutls_v._ZZN12_GLOBAL__N_110get_globalEvE6global _ZL16get_adjusted_ptrPKSt9type_infoS1_PPv _ZL21base_of_encoded_valuehP15_Unwind_Context _ZL28read_encoded_value_with_basehyPKhPy _ZL17parse_lsda_headerP15_Unwind_ContextPKhP16lsda_header_info _ZL15get_ttype_entryP16lsda_header_infoy _ZL20check_exception_specP16lsda_header_infoPKSt9type_infoPvx _ZN10__cxxabiv1L21__gxx_personality_impEiiyP17_Unwind_ExceptionP15_Unwind_Context __cxa_call_unexpected __gxx_personality_seh0 .text$_ZL16get_adjusted_ptrPKSt9type_infoS1_PPv .xdata$_ZL16get_adjusted_ptrPKSt9type_infoS1_PPv .pdata$_ZL16get_adjusted_ptrPKSt9type_infoS1_PPv .text$_ZL21base_of_encoded_valuehP15_Unwind_Context .xdata$_ZL21base_of_encoded_valuehP15_Unwind_Context .pdata$_ZL21base_C	      of_encoded_valuehP15_Unwind_Context .text$_ZL28read_encoded_value_with_basehyPKhPy .xdata$_ZL28read_encoded_value_with_basehyPKhPy .pdata$_ZL28read_encoded_value_with_basehyPKhPy .text$_ZL17parse_lsda_headerP15_Unwind_ContextPKhP16lsda_header_info .xdata$_ZL17parse_lsda_headerP15_Unwind_ContextPKhP16lsda_header_info .pdata$_ZL17parse_lsda_headerP15_Unwind_ContextPKhP16lsda_header_info .text$_ZL15get_ttype_entryP16lsda_header_infoy .xdata$_ZL15get_ttype_entryP16lsda_header_infoy .pdata$_ZL15get_ttype_entryP16lsda_header_infoy .text$_ZL20check_exception_specP16lsda_header_infoPKSt9type_infoPvx .xdata$_ZL20check_exception_specP16lsda_header_infoPKSt9type_infoPvx .pdata$_ZL20check_exception_specP16lsda_header_infoPKSt9type_infoPvx .text$_ZN10__cxxabiv1L21__gxx_personality_impEiiyP17_Unwind_ExceptionP15_Unwind_Context .xdata$_ZN10__cxxabiv1L21__gxx_personality_impEiiyP17_Unwind_ExceptionP15_Unwind_Context .pdata$_ZN10__cxxabiv1L21__gxx_personality_impEiiyP17_Unwind_ExceptionP15_Unwind_Context .text$__cxa_cD	      all_unexpected .xdata$__cxa_call_unexpected .pdata$__cxa_call_unexpected .text$__gxx_personality_seh0 .xdata$__gxx_personality_seh0 .pdata$__gxx_personality_seh0 _ZN10__cxxabiv111__terminateEPFvvE _ZSt9terminatev .rdata$.refptr._ZN10__cxxabiv119__terminate_handlerE _ZN10__cxxabiv112__unexpectedEPFvvE _ZSt10unexpectedv .rdata$.refptr._ZN10__cxxabiv120__unexpected_handlerE _ZSt13set_terminatePFvvE _ZSt13get_terminatev _ZSt14set_unexpectedPFvvE _ZSt14get_unexpectedv .text$_ZN10__cxxabiv111__terminateEPFvvE .xdata$_ZN10__cxxabiv111__terminateEPFvvE .pdata$_ZN10__cxxabiv111__terminateEPFvvE .text$_ZSt9terminatev .xdata$_ZSt9terminatev .pdata$_ZSt9terminatev .text$_ZN10__cxxabiv112__unexpectedEPFvvE .xdata$_ZN10__cxxabiv112__unexpectedEPFvvE .pdata$_ZN10__cxxabiv112__unexpectedEPFvvE .text$_ZSt10unexpectedv .xdata$_ZSt10unexpectedv .pdata$_ZSt10unexpectedv .text$_ZSt13set_terminatePFvvE .xdata$_ZSt13set_terminatePFvvE .pdata$_ZSt13set_terminatePFvvE .text$_ZSt13get_terminatev .xdata$_ZSt13get_terminatev .pdE	      ata$_ZSt13get_terminatev .text$_ZSt14set_unexpectedPFvvE .xdata$_ZSt14set_unexpectedPFvvE .pdata$_ZSt14set_unexpectedPFvvE .text$_ZSt14get_unexpectedv .xdata$_ZSt14get_unexpectedv .pdata$_ZSt14get_unexpectedv .data$_ZN10__cxxabiv119__terminate_handlerE _ZL23__gxx_exception_cleanup19_Unwind_Reason_CodeP17_Unwind_Exception __cxa_init_primary_exception __cxa_throw __cxa_rethrow .text$_ZL23__gxx_exception_cleanup19_Unwind_Reason_CodeP17_Unwind_Exception .xdata$_ZL23__gxx_exception_cleanup19_Unwind_Reason_CodeP17_Unwind_Exception .pdata$_ZL23__gxx_exception_cleanup19_Unwind_Reason_CodeP17_Unwind_Exception .text$__cxa_init_primary_exception .xdata$__cxa_init_primary_exception .pdata$__cxa_init_primary_exception .text$__cxa_throw .xdata$__cxa_throw .pdata$__cxa_throw .text$__cxa_rethrow .xdata$__cxa_rethrow .pdata$__cxa_rethrow .data$_ZN10__cxxabiv120__unexpected_handlerE .text$_ZNK9__gnu_cxx29__concurrence_broadcast_error4whatEv _ZNK9__gnu_cxx29__concurrence_broadcast_error4whatEv .text$_ZNK9__gnu_cxx24__coF	      ncurrence_wait_error4whatEv _ZNK9__gnu_cxx24__concurrence_wait_error4whatEv _ZN12_GLOBAL__N_1L4initEv _ZN12_GLOBAL__N_110fake_mutexE _ZN12_GLOBAL__N_1L12static_mutexE _ZN12_GLOBAL__N_1L16init_static_condEv _ZN12_GLOBAL__N_19fake_condE _ZN12_GLOBAL__N_1L11static_condE .text$_ZN9__gnu_cxx24__concurrence_wait_errorD1Ev _ZN9__gnu_cxx24__concurrence_wait_errorD1Ev .rdata$_ZTVN9__gnu_cxx24__concurrence_wait_errorE .text$_ZN9__gnu_cxx29__concurrence_broadcast_errorD1Ev _ZN9__gnu_cxx29__concurrence_broadcast_errorD1Ev .rdata$_ZTVN9__gnu_cxx29__concurrence_broadcast_errorE .text$_ZN9__gnu_cxx24__concurrence_wait_errorD0Ev _ZN9__gnu_cxx24__concurrence_wait_errorD0Ev .text$_ZN9__gnu_cxx29__concurrence_broadcast_errorD0Ev _ZN9__gnu_cxx29__concurrence_broadcast_errorD0Ev _ZN12_GLOBAL__N_113mutex_wrapperD2Ev.part.1 .text$_ZN9__gnu_cxx35__throw_concurrence_broadcast_errorEv _ZN9__gnu_cxx35__throw_concurrence_broadcast_errorEv .rdata$_ZTIN9__gnu_cxx29__concurrence_broadcast_errorE __cxa_guard_acquire _ZZN12_GLOBAL__NG	      _116get_static_mutexEvE4once _ZZN12_GLOBAL__N_115get_static_condEvE4once .rdata$_ZTIN9__gnu_cxx24__concurrence_wait_errorE __cxa_guard_abort __cxa_guard_release .rdata$_ZTSN9__gnu_cxx29__concurrence_broadcast_errorE .rdata$_ZTSN9__gnu_cxx24__concurrence_wait_errorE .xdata$_ZNK9__gnu_cxx29__concurrence_broadcast_error4whatEv .pdata$_ZNK9__gnu_cxx29__concurrence_broadcast_error4whatEv .xdata$_ZNK9__gnu_cxx24__concurrence_wait_error4whatEv .pdata$_ZNK9__gnu_cxx24__concurrence_wait_error4whatEv .text$_ZN12_GLOBAL__N_1L4initEv .xdata$_ZN12_GLOBAL__N_1L4initEv .pdata$_ZN12_GLOBAL__N_1L4initEv .text$_ZN12_GLOBAL__N_1L16init_static_condEv .xdata$_ZN12_GLOBAL__N_1L16init_static_condEv .pdata$_ZN12_GLOBAL__N_1L16init_static_condEv .xdata$_ZN9__gnu_cxx24__concurrence_wait_errorD1Ev .pdata$_ZN9__gnu_cxx24__concurrence_wait_errorD1Ev .xdata$_ZN9__gnu_cxx29__concurrence_broadcast_errorD1Ev .pdata$_ZN9__gnu_cxx29__concurrence_broadcast_errorD1Ev .xdata$_ZN9__gnu_cxx24__concurrence_wait_errorD0Ev .pdata$_ZN9__gnu_cxxH	      24__concurrence_wait_errorD0Ev .xdata$_ZN9__gnu_cxx29__concurrence_broadcast_errorD0Ev .pdata$_ZN9__gnu_cxx29__concurrence_broadcast_errorD0Ev .text.unlikely._ZN12_GLOBAL__N_113mutex_wrapperD2Ev.part.1 .xdata.unlikely._ZN12_GLOBAL__N_113mutex_wrapperD2Ev.part.1 .pdata.unlikely._ZN12_GLOBAL__N_113mutex_wrapperD2Ev.part.1 .xdata$_ZN9__gnu_cxx35__throw_concurrence_broadcast_errorEv .pdata$_ZN9__gnu_cxx35__throw_concurrence_broadcast_errorEv .text$__cxa_guard_acquire .xdata$__cxa_guard_acquire .pdata$__cxa_guard_acquire .text$__cxa_guard_abort .xdata$__cxa_guard_abort .pdata$__cxa_guard_abort .text$__cxa_guard_release .xdata$__cxa_guard_release .pdata$__cxa_guard_release .data$_ZZN12_GLOBAL__N_115get_static_condEvE4once .data$_ZN12_GLOBAL__N_19fake_condE .data$_ZN12_GLOBAL__N_1L11static_condE .data$_ZZN12_GLOBAL__N_116get_static_mutexEvE4once .data$_ZN12_GLOBAL__N_110fake_mutexE .data$_ZN12_GLOBAL__N_1L12static_mutexE _ZSt15set_new_handlerPFvvE _ZN12_GLOBAL__N_113__new_handlerE _ZSt15get_new_handlerv .texI	      t$_ZSt15set_new_handlerPFvvE .xdata$_ZSt15set_new_handlerPFvvE .pdata$_ZSt15set_new_handlerPFvvE .text$_ZSt15get_new_handlerv .xdata$_ZSt15get_new_handlerv .pdata$_ZSt15get_new_handlerv .data$_ZN12_GLOBAL__N_113__new_handlerE .rdata$_ZSt7nothrow .text$_Znwy .xdata$_Znwy .pdata$_Znwy .text$_Znay .xdata$_Znay .pdata$_Znay _ZnayRKSt9nothrow_t .text$_ZnayRKSt9nothrow_t .xdata$_ZnayRKSt9nothrow_t .pdata$_ZnayRKSt9nothrow_t __cxa_pure_virtual __cxa_deleted_virtual .text$__cxa_pure_virtual .xdata$__cxa_pure_virtual .pdata$__cxa_pure_virtual .text$__cxa_deleted_virtual .xdata$__cxa_deleted_virtual .pdata$__cxa_deleted_virtual _ZN10__cxxabiv120__si_class_type_infoD2Ev .rdata$_ZTVN10__cxxabiv120__si_class_type_infoE _ZN10__cxxabiv120__si_class_type_infoD1Ev _ZN10__cxxabiv120__si_class_type_infoD0Ev _ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ _ZNK10__cxxabiv120__si_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_reJ	      sultE _ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE .rdata$_ZTSN10__cxxabiv120__si_class_type_infoE .rdata$_ZTIN10__cxxabiv120__si_class_type_infoE .text$_ZN10__cxxabiv120__si_class_type_infoD2Ev .xdata$_ZN10__cxxabiv120__si_class_type_infoD2Ev .pdata$_ZN10__cxxabiv120__si_class_type_infoD2Ev .text$_ZN10__cxxabiv120__si_class_type_infoD0Ev .xdata$_ZN10__cxxabiv120__si_class_type_infoD0Ev .pdata$_ZN10__cxxabiv120__si_class_type_infoD0Ev .text$_ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .xdata$_ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .pdata$_ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .text$_ZNK10__cxxabiv120__si_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE .xdata$_ZNK10__cxxabiv120__si_class_type_info12__do_dyncastExNS_17__class_type_infK	      o10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE .pdata$_ZNK10__cxxabiv120__si_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE .text$_ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE .xdata$_ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE .pdata$_ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE _ZNSt9type_infoD2Ev _ZNSt9type_infoD1Ev _ZNKSt9type_info14__is_pointer_pEv _ZNKSt9type_info15__is_function_pEv _ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv _ZNSt9type_infoD0Ev _ZNKSt9type_infoeqERKS_ _ZNKSt9type_info10__do_catchEPKS_PPvj .rdata$_ZTVSt9type_info .text$_ZNSt9type_infoD2Ev .xdata$_ZNSt9type_infoD2Ev .pdata$_ZNSt9type_infoD2Ev .text$_ZNKSt9type_info14__is_pointer_pEv .xdata$_ZNKSt9type_info14__is_pointer_pEv .pdata$_ZNKSt9type_info14__is_pointer_pEv .textL	      $_ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .xdata$_ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .pdata$_ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .text$_ZNSt9type_infoD0Ev .xdata$_ZNSt9type_infoD0Ev .pdata$_ZNSt9type_infoD0Ev .text$_ZNKSt9type_infoeqERKS_ .xdata$_ZNKSt9type_infoeqERKS_ .pdata$_ZNKSt9type_infoeqERKS_ .text$_ZNKSt9type_info10__do_catchEPKS_PPvj .xdata$_ZNKSt9type_info10__do_catchEPKS_PPvj .pdata$_ZNKSt9type_info10__do_catchEPKS_PPvj _ZN10__cxxabiv121__vmi_class_type_infoD2Ev .rdata$_ZTVN10__cxxabiv121__vmi_class_type_infoE _ZN10__cxxabiv121__vmi_class_type_infoD1Ev _ZN10__cxxabiv121__vmi_class_type_infoD0Ev _ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ _ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE _ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_1M	      6__dyncast_resultE .rdata$_ZTSN10__cxxabiv121__vmi_class_type_infoE .rdata$_ZTIN10__cxxabiv121__vmi_class_type_infoE .text$_ZN10__cxxabiv121__vmi_class_type_infoD2Ev .xdata$_ZN10__cxxabiv121__vmi_class_type_infoD2Ev .pdata$_ZN10__cxxabiv121__vmi_class_type_infoD2Ev .text$_ZN10__cxxabiv121__vmi_class_type_infoD0Ev .xdata$_ZN10__cxxabiv121__vmi_class_type_infoD0Ev .pdata$_ZN10__cxxabiv121__vmi_class_type_infoD0Ev .text$_ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .xdata$_ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .pdata$_ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcExPKvPKNS_17__class_type_infoES2_ .text$_ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE .xdata$_ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE .pdata$_ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__clasN	      s_type_infoEPKvRNS1_15__upcast_resultE .text$_ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE .xdata$_ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE .pdata$_ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastExNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE _ZN9__gnu_cxx27__verbose_terminate_handlerEv _ZZN9__gnu_cxx27__verbose_terminate_handlerEvE11terminating .text$_ZN9__gnu_cxx27__verbose_terminate_handlerEv .xdata$_ZN9__gnu_cxx27__verbose_terminate_handlerEv .pdata$_ZN9__gnu_cxx27__verbose_terminate_handlerEv .data$_ZZN9__gnu_cxx27__verbose_terminate_handlerEvE11terminating _ZN12_GLOBAL__N_1L10fopen_modeESt13_Ios_Openmode _ZN12_GLOBAL__N_1L6xwriteEiPKcx _ZNSt12__basic_fileIcEC2EPPv _ZNSt12__basic_fileIcEC1EPPv _ZNSt12__basic_fileIcE8sys_openEP6_iobufSt13_Ios_Openmode _ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_OpenmO	      ode _ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei _ZNKSt12__basic_fileIcE7is_openEv _ZNSt12__basic_fileIcE2fdEv _ZNSt12__basic_fileIcE4fileEv _ZNSt12__basic_fileIcE5closeEv _ZNSt12__basic_fileIcED2Ev _ZNSt12__basic_fileIcED1Ev _ZNSt12__basic_fileIcE6xsgetnEPcx _ZNSt12__basic_fileIcE6xsputnEPKcx _ZNSt12__basic_fileIcE8xsputn_2EPKcxS2_x _ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir _ZNSt12__basic_fileIcE4syncEv _ZNSt12__basic_fileIcE9showmanycEv .text$_ZN12_GLOBAL__N_1L10fopen_modeESt13_Ios_Openmode .xdata$_ZN12_GLOBAL__N_1L10fopen_modeESt13_Ios_Openmode .pdata$_ZN12_GLOBAL__N_1L10fopen_modeESt13_Ios_Openmode .text$_ZN12_GLOBAL__N_1L6xwriteEiPKcx .xdata$_ZN12_GLOBAL__N_1L6xwriteEiPKcx .pdata$_ZN12_GLOBAL__N_1L6xwriteEiPKcx .text$_ZNSt12__basic_fileIcEC2EPPv .xdata$_ZNSt12__basic_fileIcEC2EPPv .pdata$_ZNSt12__basic_fileIcEC2EPPv .text$_ZNSt12__basic_fileIcE8sys_openEP6_iobufSt13_Ios_Openmode .xdata$_ZNSt12__basic_fileIcE8sys_openEP6_iobufSt13_Ios_Openmode .pdata$_ZNSt12__basic_fileIcE8sys_openEP6_P	      iobufSt13_Ios_Openmode .text$_ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_Openmode .xdata$_ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_Openmode .pdata$_ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_Openmode .text$_ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei .xdata$_ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei .pdata$_ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei .text$_ZNKSt12__basic_fileIcE7is_openEv .xdata$_ZNKSt12__basic_fileIcE7is_openEv .pdata$_ZNKSt12__basic_fileIcE7is_openEv .text$_ZNSt12__basic_fileIcE2fdEv .xdata$_ZNSt12__basic_fileIcE2fdEv .pdata$_ZNSt12__basic_fileIcE2fdEv .text$_ZNSt12__basic_fileIcE4fileEv .xdata$_ZNSt12__basic_fileIcE4fileEv .pdata$_ZNSt12__basic_fileIcE4fileEv .text$_ZNSt12__basic_fileIcE5closeEv .xdata$_ZNSt12__basic_fileIcE5closeEv .pdata$_ZNSt12__basic_fileIcE5closeEv .text$_ZNSt12__basic_fileIcED2Ev .xdata$_ZNSt12__basic_fileIcED2Ev .pdata$_ZNSt12__basic_fileIcED2Ev .text$_ZNSt12__basic_fileIcE6xsgetnEPcx .xdata$_ZNSt12__basic_fileIcE6xsgetnEPcx .pdata$_ZNSt12__basQ	      ic_fileIcE6xsgetnEPcx .text$_ZNSt12__basic_fileIcE6xsputnEPKcx .xdata$_ZNSt12__basic_fileIcE6xsputnEPKcx .pdata$_ZNSt12__basic_fileIcE6xsputnEPKcx .text$_ZNSt12__basic_fileIcE8xsputn_2EPKcxS2_x .xdata$_ZNSt12__basic_fileIcE8xsputn_2EPKcxS2_x .pdata$_ZNSt12__basic_fileIcE8xsputn_2EPKcxS2_x .text$_ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir .xdata$_ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir .pdata$_ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir .text$_ZNSt12__basic_fileIcE4syncEv .xdata$_ZNSt12__basic_fileIcE4syncEv .pdata$_ZNSt12__basic_fileIcE4syncEv .text$_ZNSt12__basic_fileIcE9showmanycEv .xdata$_ZNSt12__basic_fileIcE9showmanycEv .pdata$_ZNSt12__basic_fileIcE9showmanycEv _ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi _ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi _ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi _ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ _ZNSt6locale5facet19_S_destroy_c_localeERPi _ZNSt6locale5facet17_S_clone_c_localeERPi _ZNSt6locale5facet20_S_lc_ctype_cR	      _localeEPiPKc _ZN9__gnu_cxxL14category_namesE .text$_ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi .xdata$_ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi .pdata$_ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi .text$_ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi .xdata$_ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi .pdata$_ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi .text$_ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi .xdata$_ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi .pdata$_ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi .text$_ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ .xdata$_ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ .pdata$_ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ .text$_ZNSt6locale5facet19_S_destroy_c_localeERPi .xdata$_ZNSt6locale5facet19_S_destroy_c_localeERPi .pdata$_ZNSt6locale5facet19_S_destroy_c_localeERPi .text$_ZNSt6locale5facet17_S_clone_c_localeERPi .xdata$_ZNSt6locale5facet17_S_clone_c_localeERPi .pdata$_ZNSt6locale5facet1S	      7_S_clone_c_localeERPi .text$_ZNSt6locale5facet20_S_lc_ctype_c_localeEPiPKc .xdata$_ZNSt6locale5facet20_S_lc_ctype_c_localeEPiPKc .pdata$_ZNSt6locale5facet20_S_lc_ctype_c_localeEPiPKc .rdata$_ZNSt6locale13_S_categoriesE .rdata$_ZN9__gnu_cxxL14category_namesE _ZNKSt7codecvtIcciE6do_outERiPKcS3_RS3_PcS5_RS5_ _ZNKSt7codecvtIcciE5do_inERiPKcS3_RS3_PcS5_RS5_ _ZNKSt7codecvtIcciE10do_unshiftERiPcS2_RS2_ _ZNKSt7codecvtIwciE10do_unshiftERiPcS2_RS2_ _ZNKSt7codecvtIcciE11do_encodingEv _ZNKSt7codecvtIcciE13do_max_lengthEv _ZNKSt7codecvtIcciE16do_always_noconvEv _ZNKSt7codecvtIcciE9do_lengthERiPKcS3_y _ZNKSt7codecvtIwciE16do_always_noconvEv _ZNSt7codecvtIcciED2Ev .rdata$_ZTVSt7codecvtIcciE .rdata$.refptr._ZTVSt23__codecvt_abstract_baseIcciE _ZNSt7codecvtIcciED1Ev _ZNSt7codecvtIwciED2Ev .rdata$_ZTVSt7codecvtIwciE .rdata$.refptr._ZTVSt23__codecvt_abstract_baseIwciE _ZNSt7codecvtIwciED1Ev _ZNSt7codecvtIcciED0Ev _ZNSt7codecvtIwciED0Ev _ZNSt7codecvtIcciEC2Ey _ZNSt7codecvtIcciEC1Ey _ZNSt7codecvtIcciEC2EPiy _ZNSt7codecvtT	      IcciEC1EPiy _ZNSt7codecvtIwciEC2Ey _ZNSt7codecvtIwciEC1Ey _ZNSt7codecvtIwciEC2EPiy _ZNSt7codecvtIwciEC1EPiy .text$_ZNKSt7codecvtIcciE6do_outERiPKcS3_RS3_PcS5_RS5_ .xdata$_ZNKSt7codecvtIcciE6do_outERiPKcS3_RS3_PcS5_RS5_ .pdata$_ZNKSt7codecvtIcciE6do_outERiPKcS3_RS3_PcS5_RS5_ .text$_ZNKSt7codecvtIcciE10do_unshiftERiPcS2_RS2_ .xdata$_ZNKSt7codecvtIcciE10do_unshiftERiPcS2_RS2_ .pdata$_ZNKSt7codecvtIcciE10do_unshiftERiPcS2_RS2_ .text$_ZNKSt7codecvtIcciE11do_encodingEv .xdata$_ZNKSt7codecvtIcciE11do_encodingEv .pdata$_ZNKSt7codecvtIcciE11do_encodingEv .text$_ZNKSt7codecvtIcciE16do_always_noconvEv .xdata$_ZNKSt7codecvtIcciE16do_always_noconvEv .pdata$_ZNKSt7codecvtIcciE16do_always_noconvEv .text$_ZNKSt7codecvtIcciE9do_lengthERiPKcS3_y .xdata$_ZNKSt7codecvtIcciE9do_lengthERiPKcS3_y .pdata$_ZNKSt7codecvtIcciE9do_lengthERiPKcS3_y .text$_ZNKSt7codecvtIwciE16do_always_noconvEv .xdata$_ZNKSt7codecvtIwciE16do_always_noconvEv .pdata$_ZNKSt7codecvtIwciE16do_always_noconvEv .text$_ZNSt7codecvtIcciED2Ev .xdata$_ZNSt7coU	      decvtIcciED2Ev .pdata$_ZNSt7codecvtIcciED2Ev .text$_ZNSt7codecvtIwciED2Ev .xdata$_ZNSt7codecvtIwciED2Ev .pdata$_ZNSt7codecvtIwciED2Ev .text$_ZNSt7codecvtIcciED0Ev .xdata$_ZNSt7codecvtIcciED0Ev .pdata$_ZNSt7codecvtIcciED0Ev .text$_ZNSt7codecvtIwciED0Ev .xdata$_ZNSt7codecvtIwciED0Ev .pdata$_ZNSt7codecvtIwciED0Ev .text$_ZNSt7codecvtIcciEC2Ey .xdata$_ZNSt7codecvtIcciEC2Ey .pdata$_ZNSt7codecvtIcciEC2Ey .text$_ZNSt7codecvtIcciEC2EPiy .xdata$_ZNSt7codecvtIcciEC2EPiy .pdata$_ZNSt7codecvtIcciEC2EPiy .text$_ZNSt7codecvtIwciEC2Ey .xdata$_ZNSt7codecvtIwciEC2Ey .pdata$_ZNSt7codecvtIwciEC2Ey .text$_ZNSt7codecvtIwciEC2EPiy .xdata$_ZNSt7codecvtIwciEC2EPiy .pdata$_ZNSt7codecvtIwciEC2EPiy .data$_ZNSt7codecvtIwciE2idE .data$_ZNSt7codecvtIcciE2idE _ZNKSt7codecvtIwciE6do_outERiPKwS3_RS3_PcS5_RS5_ _ZNKSt7codecvtIwciE5do_inERiPKcS3_RS3_PwS5_RS5_ _ZNKSt7codecvtIwciE11do_encodingEv _ZNKSt7codecvtIwciE13do_max_lengthEv _ZNKSt7codecvtIwciE9do_lengthERiPKcS3_y .text$_ZNKSt7codecvtIwciE6do_outERiPKwS3_RS3_PcS5_RS5_ .xdata$_ZNKSt7V	      codecvtIwciE6do_outERiPKwS3_RS3_PcS5_RS5_ .pdata$_ZNKSt7codecvtIwciE6do_outERiPKwS3_RS3_PcS5_RS5_ .text$_ZNKSt7codecvtIwciE5do_inERiPKcS3_RS3_PwS5_RS5_ .xdata$_ZNKSt7codecvtIwciE5do_inERiPKcS3_RS3_PwS5_RS5_ .pdata$_ZNKSt7codecvtIwciE5do_inERiPKcS3_RS3_PwS5_RS5_ .text$_ZNKSt7codecvtIwciE11do_encodingEv .xdata$_ZNKSt7codecvtIwciE11do_encodingEv .pdata$_ZNKSt7codecvtIwciE11do_encodingEv .text$_ZNKSt7codecvtIwciE13do_max_lengthEv .xdata$_ZNKSt7codecvtIwciE13do_max_lengthEv .pdata$_ZNKSt7codecvtIwciE13do_max_lengthEv .text$_ZNKSt7codecvtIwciE9do_lengthERiPKcS3_y .xdata$_ZNKSt7codecvtIwciE9do_lengthERiPKcS3_y .pdata$_ZNKSt7codecvtIwciE9do_lengthERiPKcS3_y _ZNKSt7__cxx117collateIcE10_M_compareEPKcS3_ _ZNKSt7__cxx117collateIcE12_M_transformEPcPKcy _ZNKSt7__cxx117collateIwE10_M_compareEPKwS3_ _ZNKSt7__cxx117collateIwE12_M_transformEPwPKwy .text$_ZNKSt7__cxx117collateIcE10_M_compareEPKcS3_ .xdata$_ZNKSt7__cxx117collateIcE10_M_compareEPKcS3_ .pdata$_ZNKSt7__cxx117collateIcE10_M_compareEPKcS3_ .text$_ZNKSt7__cxx1W	      17collateIcE12_M_transformEPcPKcy .xdata$_ZNKSt7__cxx117collateIcE12_M_transformEPcPKcy .pdata$_ZNKSt7__cxx117collateIcE12_M_transformEPcPKcy .text$_ZNKSt7__cxx117collateIwE10_M_compareEPKwS3_ .xdata$_ZNKSt7__cxx117collateIwE10_M_compareEPKwS3_ .pdata$_ZNKSt7__cxx117collateIwE10_M_compareEPKwS3_ .text$_ZNKSt7__cxx117collateIwE12_M_transformEPwPKwy .xdata$_ZNKSt7__cxx117collateIwE12_M_transformEPwPKwy .pdata$_ZNKSt7__cxx117collateIwE12_M_transformEPwPKwy _ZNKSt7collateIcE10_M_compareEPKcS2_ _ZNKSt7collateIcE12_M_transformEPcPKcy _ZNKSt7collateIwE10_M_compareEPKwS2_ _ZNKSt7collateIwE12_M_transformEPwPKwy .text$_ZNKSt7collateIcE10_M_compareEPKcS2_ .xdata$_ZNKSt7collateIcE10_M_compareEPKcS2_ .pdata$_ZNKSt7collateIcE10_M_compareEPKcS2_ .text$_ZNKSt7collateIcE12_M_transformEPcPKcy .xdata$_ZNKSt7collateIcE12_M_transformEPcPKcy .pdata$_ZNKSt7collateIcE12_M_transformEPcPKcy .text$_ZNKSt7collateIwE10_M_compareEPKwS2_ .xdata$_ZNKSt7collateIwE10_M_compareEPKwS2_ .pdata$_ZNKSt7collateIwE10_M_compareEPKwS2_ .text$_X	      ZNKSt7collateIwE12_M_transformEPwPKwy .xdata$_ZNKSt7collateIwE12_M_transformEPwPKwy .pdata$_ZNKSt7collateIwE12_M_transformEPwPKwy _ZNSt8ios_base7_M_initEv _ZNSt8ios_base5imbueERKSt6locale .text$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv _ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv .text$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvPvEv _ZNKSt9basic_iosIwSt11char_traitsIwEEcvPvEv .text$_ZNSt8ios_base7_M_initEv .xdata$_ZNSt8ios_base7_M_initEv .pdata$_ZNSt8ios_base7_M_initEv .text$_ZNSt8ios_base5imbueERKSt6locale .xdata$_ZNSt8ios_base5imbueERKSt6locale .pdata$_ZNSt8ios_base5imbueERKSt6locale .xdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv .pdata$_ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv .xdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvPvEv .pdata$_ZNKSt9basic_iosIwSt11char_traitsIwEEcvPvEv _ZNSi7getlineEPcxc _ZNSi6ignoreExi _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ _ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwxw _ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreExt .text$_ZNSi7getlineEY	      Pcxc .xdata$_ZNSi7getlineEPcxc .pdata$_ZNSi7getlineEPcxc .text$_ZNSi6ignoreExi .xdata$_ZNSi6ignoreExi .pdata$_ZNSi6ignoreExi .text$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ .xdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ .pdata$_ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwxw .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwxw .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE7getlineEPwxw .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreExt .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreExt .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreExt _ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc _ZSt22__verify_grouping_implPKcyS0_y _ZSt17__verify_groupingPKcyRKSs .text$_ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc .xdata$_ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc .pdata$_ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc .text$_ZSt22__verify_grouping_impZ	      lPKcyS0_y .xdata$_ZSt22__verify_grouping_implPKcyS0_y .pdata$_ZSt22__verify_grouping_implPKcyS0_y .text$_ZSt17__verify_groupingPKcyRKSs .xdata$_ZSt17__verify_groupingPKcyRKSs .pdata$_ZSt17__verify_groupingPKcyRKSs .data$_ZNSt10__num_base12_S_atoms_outE .data$_ZNSt10__num_base11_S_atoms_inE .data$_ZNSt10money_base8_S_atomsE .rdata$_ZNSt10money_base18_S_default_patternE .data$_ZNSt17__timepunct_cacheIwE12_S_timezonesE .data$_ZNSt17__timepunct_cacheIcE12_S_timezonesE _ZNKSt7__cxx118messagesIcE6do_getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE _ZNKSt7__cxx118messagesIwE6do_getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .text$_ZNKSt7__cxx118messagesIcE6do_getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNKSt7__cxx118messagesIcE6do_getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNKSt7__cxx118messagesIcE6do_getEiiiRKNS_12basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNKSt7__cxx118messagesIwE6do_getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .xdata$_ZNKSt7__c[	      xx118messagesIwE6do_getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE .pdata$_ZNKSt7__cxx118messagesIwE6do_getEiiiRKNS_12basic_stringIwSt11char_traitsIwESaIwEEE _ZNKSt8messagesIcE6do_getEiiiRKSs _ZNKSt8messagesIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .text$_ZNKSt8messagesIcE6do_getEiiiRKSs .xdata$_ZNKSt8messagesIcE6do_getEiiiRKSs .pdata$_ZNKSt8messagesIcE6do_getEiiiRKSs .text$_ZNKSt8messagesIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .xdata$_ZNKSt8messagesIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .pdata$_ZNKSt8messagesIwE6do_getEiiiRKSbIwSt11char_traitsIwESaIwEE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EE .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_ .text$_ZNSt7__cxx1112\	      basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEyc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEyc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvS9_T_SA_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvS9_T_SA_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_RKS4_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_RKS4_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcy _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE]	      7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcy .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_yc _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_yc .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S7_S7_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S7_S7_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcSA_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcSA_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9_^	      _gnu_cxx17__normal_iteratorIPcS4_EES8_S8_S8_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S8_S8_ .text$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_NS6_IPKcS4_EESB_ _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_NS6_IPKcS4_EESB_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EE .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEyw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIP_	      wS4_EEyw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvS9_T_SA_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvS9_T_SA_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_RKS4_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_RKS4_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwy _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwy .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKw _ZNSt7__cxx1`	      112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_yw _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_yw .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S7_S7_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S7_S7_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwSA_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwSA_ .text$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S8_S8_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S8_S8_ .text$_ZNSt7__cxx1112basia	      c_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_NS6_IPKwS4_EESB_ _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_NS6_IPKwS4_EESB_ _ZSt17__verify_groupingPKcyRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EE .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EE .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE5eraseEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEyc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEyc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6inseb	      rtIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvS9_T_SA_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertIN9__gnu_cxx17__normal_iteratorIPcS4_EEEEvS9_T_SA_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE6insertEN9__gnu_cxx17__normal_iteratorIPcS4_EEc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_RKS4_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_RKS4_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcy .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcy .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcc	      ESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_yc .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_yc .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S7_S7_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S7_S7_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcSA_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_PKcSA_ .xdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S8_S8_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_S8_S8_ .xdata$_ZNSt7__cxx1112basicd	      _stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_NS6_IPKcS4_EESB_ .pdata$_ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE7replaceEN9__gnu_cxx17__normal_iteratorIPcS4_EES8_NS6_IPKcS4_EESB_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EE .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EE .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE5eraseEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEyw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEyw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvS9_T_SA_ .pdata$_ZNSt7__cxx1112be	      asic_stringIwSt11char_traitsIwESaIwEE6insertIN9__gnu_cxx17__normal_iteratorIPwS4_EEEEvS9_T_SA_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE6insertEN9__gnu_cxx17__normal_iteratorIPwS4_EEw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_RKS4_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_RKS4_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwy .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwy .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKw .xdata$_ZNSt7__f	      cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_yw .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_yw .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S7_S7_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S7_S7_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwSA_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_PKwSA_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S8_S8_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_S8_S8_ .xdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwSg	      4_EES8_NS6_IPKwS4_EESB_ .pdata$_ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE7replaceEN9__gnu_cxx17__normal_iteratorIPwS4_EES8_NS6_IPKwS4_EESB_ .text$_ZSt17__verify_groupingPKcyRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZSt17__verify_groupingPKcyRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZSt17__verify_groupingPKcyRKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNKSt11logic_error4whatEv _ZNKSt13runtime_error4whatEv _ZNSt11logic_errorD2Ev .rdata$_ZTVSt11logic_error _ZNSt11logic_errorD1Ev _ZNSt12domain_errorD2Ev .rdata$_ZTVSt12domain_error _ZNSt12domain_errorD1Ev _ZNSt16invalid_argumentD2Ev .rdata$_ZTVSt16invalid_argument _ZNSt16invalid_argumentD1Ev _ZNSt12length_errorD2Ev .rdata$_ZTVSt12length_error _ZNSt12length_errorD1Ev _ZNSt12out_of_rangeD2Ev .rdata$_ZTVSt12out_of_range _ZNSt12out_of_rangeD1Ev _ZNSt11logic_errorD0Ev _ZNSt12domain_errorD0Ev _ZNSt16invalid_argumentD0Ev _ZNSt12length_errorD0Ev _ZNSt12out_of_rangeD0Ev _ZNSt13runtime_errorD2Ev .rdatah	      $_ZTVSt13runtime_error _ZNSt13runtime_errorD1Ev _ZNSt13runtime_errorD0Ev _ZNSt11range_errorD2Ev .rdata$_ZTVSt11range_error _ZNSt11range_errorD1Ev _ZNSt11range_errorD0Ev _ZNSt14overflow_errorD2Ev .rdata$_ZTVSt14overflow_error _ZNSt14overflow_errorD1Ev _ZNSt14overflow_errorD0Ev _ZNSt15underflow_errorD2Ev .rdata$_ZTVSt15underflow_error _ZNSt15underflow_errorD1Ev _ZNSt15underflow_errorD0Ev _ZNSt11logic_errorC2ERKSs _ZNSt11logic_errorC1ERKSs _ZNSt12domain_errorC2ERKSs _ZNSt12domain_errorC1ERKSs _ZNSt16invalid_argumentC2ERKSs _ZNSt16invalid_argumentC1ERKSs _ZNSt12length_errorC2ERKSs _ZNSt12length_errorC1ERKSs _ZNSt12out_of_rangeC2ERKSs _ZNSt12out_of_rangeC1ERKSs _ZNSt13runtime_errorC2ERKSs _ZNSt13runtime_errorC1ERKSs _ZNSt11range_errorC2ERKSs _ZNSt11range_errorC1ERKSs _ZNSt14overflow_errorC2ERKSs _ZNSt14overflow_errorC1ERKSs _ZNSt15underflow_errorC2ERKSs _ZNSt15underflow_errorC1ERKSs .text$_ZNKSt11logic_error4whatEv .xdata$_ZNKSt11logic_error4whatEv .pdata$_ZNKSt11logic_error4whatEv .text$_ZNKSt13runtime_eri	      ror4whatEv .xdata$_ZNKSt13runtime_error4whatEv .pdata$_ZNKSt13runtime_error4whatEv .text$_ZNSt11logic_errorD2Ev .xdata$_ZNSt11logic_errorD2Ev .pdata$_ZNSt11logic_errorD2Ev .text$_ZNSt12domain_errorD2Ev .xdata$_ZNSt12domain_errorD2Ev .pdata$_ZNSt12domain_errorD2Ev .text$_ZNSt16invalid_argumentD2Ev .xdata$_ZNSt16invalid_argumentD2Ev .pdata$_ZNSt16invalid_argumentD2Ev .text$_ZNSt12length_errorD2Ev .xdata$_ZNSt12length_errorD2Ev .pdata$_ZNSt12length_errorD2Ev .text$_ZNSt12out_of_rangeD2Ev .xdata$_ZNSt12out_of_rangeD2Ev .pdata$_ZNSt12out_of_rangeD2Ev .text$_ZNSt11logic_errorD0Ev .xdata$_ZNSt11logic_errorD0Ev .pdata$_ZNSt11logic_errorD0Ev .text$_ZNSt12domain_errorD0Ev .xdata$_ZNSt12domain_errorD0Ev .pdata$_ZNSt12domain_errorD0Ev .text$_ZNSt16invalid_argumentD0Ev .xdata$_ZNSt16invalid_argumentD0Ev .pdata$_ZNSt16invalid_argumentD0Ev .text$_ZNSt12length_errorD0Ev .xdata$_ZNSt12length_errorD0Ev .pdata$_ZNSt12length_errorD0Ev .text$_ZNSt12out_of_rangeD0Ev .xdata$_ZNSt12out_of_rangeD0Ev .pdata$_ZNSt12out_of_rangej	      D0Ev .text$_ZNSt13runtime_errorD2Ev .xdata$_ZNSt13runtime_errorD2Ev .pdata$_ZNSt13runtime_errorD2Ev .text$_ZNSt13runtime_errorD0Ev .xdata$_ZNSt13runtime_errorD0Ev .pdata$_ZNSt13runtime_errorD0Ev .text$_ZNSt11range_errorD2Ev .xdata$_ZNSt11range_errorD2Ev .pdata$_ZNSt11range_errorD2Ev .text$_ZNSt11range_errorD0Ev .xdata$_ZNSt11range_errorD0Ev .pdata$_ZNSt11range_errorD0Ev .text$_ZNSt14overflow_errorD2Ev .xdata$_ZNSt14overflow_errorD2Ev .pdata$_ZNSt14overflow_errorD2Ev .text$_ZNSt14overflow_errorD0Ev .xdata$_ZNSt14overflow_errorD0Ev .pdata$_ZNSt14overflow_errorD0Ev .text$_ZNSt15underflow_errorD2Ev .xdata$_ZNSt15underflow_errorD2Ev .pdata$_ZNSt15underflow_errorD2Ev .text$_ZNSt15underflow_errorD0Ev .xdata$_ZNSt15underflow_errorD0Ev .pdata$_ZNSt15underflow_errorD0Ev .text$_ZNSt11logic_errorC2ERKSs .xdata$_ZNSt11logic_errorC2ERKSs .pdata$_ZNSt11logic_errorC2ERKSs .text$_ZNSt12domain_errorC2ERKSs .xdata$_ZNSt12domain_errorC2ERKSs .pdata$_ZNSt12domain_errorC2ERKSs .text$_ZNSt16invalid_argumentC2ERKSs .xdata$_Zk	      NSt16invalid_argumentC2ERKSs .pdata$_ZNSt16invalid_argumentC2ERKSs .text$_ZNSt12length_errorC2ERKSs .xdata$_ZNSt12length_errorC2ERKSs .pdata$_ZNSt12length_errorC2ERKSs .text$_ZNSt12out_of_rangeC2ERKSs .xdata$_ZNSt12out_of_rangeC2ERKSs .pdata$_ZNSt12out_of_rangeC2ERKSs .text$_ZNSt13runtime_errorC2ERKSs .xdata$_ZNSt13runtime_errorC2ERKSs .pdata$_ZNSt13runtime_errorC2ERKSs .text$_ZNSt11range_errorC2ERKSs .xdata$_ZNSt11range_errorC2ERKSs .pdata$_ZNSt11range_errorC2ERKSs .text$_ZNSt14overflow_errorC2ERKSs .xdata$_ZNSt14overflow_errorC2ERKSs .pdata$_ZNSt14overflow_errorC2ERKSs .text$_ZNSt15underflow_errorC2ERKSs .xdata$_ZNSt15underflow_errorC2ERKSs .pdata$_ZNSt15underflow_errorC2ERKSs _ZSt21__copy_streambufs_eofIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_Rb _ZSt21__copy_streambufs_eofIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_Rb .text$_ZSt21__copy_streambufs_eofIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_Rb .xdata$_ZSt21__copy_streambufs_eofIcSt11char_traitsIcEExPSt15basic_streambufl	      IT_T0_ES6_Rb .pdata$_ZSt21__copy_streambufs_eofIcSt11char_traitsIcEExPSt15basic_streambufIT_T0_ES6_Rb .text$_ZSt21__copy_streambufs_eofIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_Rb .xdata$_ZSt21__copy_streambufs_eofIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_Rb .pdata$_ZSt21__copy_streambufs_eofIwSt11char_traitsIwEExPSt15basic_streambufIT_T0_ES6_Rb _ZNKSt11__timepunctIcE6_M_putEPcyPKcPK2tm _ZNSt11__timepunctIcE23_M_initialize_timepunctEPi _ZNKSt11__timepunctIwE6_M_putEPwyPKwPK2tm _ZNSt11__timepunctIwE23_M_initialize_timepunctEPi .text$_ZNKSt11__timepunctIcE6_M_putEPcyPKcPK2tm .xdata$_ZNKSt11__timepunctIcE6_M_putEPcyPKcPK2tm .pdata$_ZNKSt11__timepunctIcE6_M_putEPcyPKcPK2tm .text$_ZNSt11__timepunctIcE23_M_initialize_timepunctEPi .xdata$_ZNSt11__timepunctIcE23_M_initialize_timepunctEPi .pdata$_ZNSt11__timepunctIcE23_M_initialize_timepunctEPi .text$_ZNKSt11__timepunctIwE6_M_putEPwyPKwPK2tm .xdata$_ZNKSt11__timepunctIwE6_M_putEPwyPKwPK2tm .pdata$_ZNKSt11__timepunctIwE6_M_putEPwyPKwPK2tm .tm	      ext$_ZNSt11__timepunctIwE23_M_initialize_timepunctEPi .xdata$_ZNSt11__timepunctIwE23_M_initialize_timepunctEPi .pdata$_ZNSt11__timepunctIwE23_M_initialize_timepunctEPi _ZNSt11logic_errorC2ERKS_ .rdata$.refptr._ZTVSt11logic_error _ZNSt11logic_errorC1ERKS_ _ZNSt11logic_erroraSERKS_ _ZNSt13runtime_errorC2ERKS_ .rdata$.refptr._ZTVSt13runtime_error _ZNSt13runtime_errorC1ERKS_ _ZNSt13runtime_erroraSERKS_ _ZNSt11logic_errorC2EPKc _ZNSt11logic_errorC1EPKc _ZNSt12domain_errorC2EPKc .rdata$.refptr._ZTVSt12domain_error _ZNSt12domain_errorC1EPKc _ZNSt16invalid_argumentC2EPKc .rdata$.refptr._ZTVSt16invalid_argument _ZNSt16invalid_argumentC1EPKc _ZNSt12length_errorC2EPKc .rdata$.refptr._ZTVSt12length_error _ZNSt12length_errorC1EPKc _ZNSt12out_of_rangeC2EPKc .rdata$.refptr._ZTVSt12out_of_range _ZNSt12out_of_rangeC1EPKc _ZNSt13runtime_errorC2EPKc _ZNSt13runtime_errorC1EPKc _ZNSt11range_errorC2EPKc .rdata$.refptr._ZTVSt11range_error _ZNSt11range_errorC1EPKc _ZNSt14overflow_errorC2EPKc .rdata$.refptr._ZTVSt14overflow_en	      rror _ZNSt14overflow_errorC1EPKc _ZNSt15underflow_errorC2EPKc .rdata$.refptr._ZTVSt15underflow_error _ZNSt15underflow_errorC1EPKc _ZNSt12__sso_stringC2ERKSs _ZNSt12__sso_stringC1ERKSs _ZNSt12__cow_stringC2Ev _ZNSt12__cow_stringC1Ev _ZNSt12__cow_stringC2ERKSs _ZNSt12__cow_stringC1ERKSs _ZNSt12__cow_stringC2EPKcy _ZNSt12__cow_stringC1EPKcy _ZNSt12__cow_stringC2ERKS_ _ZNSt12__cow_stringC1ERKS_ _ZNSt12__cow_stringaSERKS_ _ZNSt12__cow_stringD2Ev _ZNSt12__cow_stringD1Ev _ZNSt12__cow_stringC2EOS_ _ZNSt12__cow_stringC1EOS_ _ZNSt12__cow_stringaSEOS_ _ZNKSt3_V214error_category10_M_messageEi .text$_ZNSt11logic_errorC2ERKS_ .xdata$_ZNSt11logic_errorC2ERKS_ .pdata$_ZNSt11logic_errorC2ERKS_ .text$_ZNSt11logic_erroraSERKS_ .xdata$_ZNSt11logic_erroraSERKS_ .pdata$_ZNSt11logic_erroraSERKS_ .text$_ZNSt13runtime_errorC2ERKS_ .xdata$_ZNSt13runtime_errorC2ERKS_ .pdata$_ZNSt13runtime_errorC2ERKS_ .text$_ZNSt13runtime_erroraSERKS_ .xdata$_ZNSt13runtime_erroraSERKS_ .pdata$_ZNSt13runtime_erroraSERKS_ .text$_ZNSt11logic_erroro	      C2EPKc .xdata$_ZNSt11logic_errorC2EPKc .pdata$_ZNSt11logic_errorC2EPKc .text$_ZNSt12domain_errorC2EPKc .xdata$_ZNSt12domain_errorC2EPKc .pdata$_ZNSt12domain_errorC2EPKc .text$_ZNSt16invalid_argumentC2EPKc .xdata$_ZNSt16invalid_argumentC2EPKc .pdata$_ZNSt16invalid_argumentC2EPKc .text$_ZNSt12length_errorC2EPKc .xdata$_ZNSt12length_errorC2EPKc .pdata$_ZNSt12length_errorC2EPKc .text$_ZNSt12out_of_rangeC2EPKc .xdata$_ZNSt12out_of_rangeC2EPKc .pdata$_ZNSt12out_of_rangeC2EPKc .text$_ZNSt13runtime_errorC2EPKc .xdata$_ZNSt13runtime_errorC2EPKc .pdata$_ZNSt13runtime_errorC2EPKc .text$_ZNSt11range_errorC2EPKc .xdata$_ZNSt11range_errorC2EPKc .pdata$_ZNSt11range_errorC2EPKc .text$_ZNSt14overflow_errorC2EPKc .xdata$_ZNSt14overflow_errorC2EPKc .pdata$_ZNSt14overflow_errorC2EPKc .text$_ZNSt15underflow_errorC2EPKc .xdata$_ZNSt15underflow_errorC2EPKc .pdata$_ZNSt15underflow_errorC2EPKc .text$_ZNSt12__sso_stringC2ERKSs .xdata$_ZNSt12__sso_stringC2ERKSs .pdata$_ZNSt12__sso_stringC2ERKSs .text$_ZNSt12__cow_stringC2Ev .xdp	      ata$_ZNSt12__cow_stringC2Ev .pdata$_ZNSt12__cow_stringC2Ev .text$_ZNSt12__cow_stringC2ERKSs .xdata$_ZNSt12__cow_stringC2ERKSs .pdata$_ZNSt12__cow_stringC2ERKSs .text$_ZNSt12__cow_stringC2EPKcy .xdata$_ZNSt12__cow_stringC2EPKcy .pdata$_ZNSt12__cow_stringC2EPKcy .text$_ZNSt12__cow_stringC2ERKS_ .xdata$_ZNSt12__cow_stringC2ERKS_ .pdata$_ZNSt12__cow_stringC2ERKS_ .text$_ZNSt12__cow_stringaSERKS_ .xdata$_ZNSt12__cow_stringaSERKS_ .pdata$_ZNSt12__cow_stringaSERKS_ .text$_ZNSt12__cow_stringD2Ev .xdata$_ZNSt12__cow_stringD2Ev .pdata$_ZNSt12__cow_stringD2Ev .text$_ZNSt12__cow_stringC2EOS_ .xdata$_ZNSt12__cow_stringC2EOS_ .pdata$_ZNSt12__cow_stringC2EOS_ .text$_ZNSt12__cow_stringaSEOS_ .xdata$_ZNSt12__cow_stringaSEOS_ .pdata$_ZNSt12__cow_stringaSEOS_ .text$_ZNKSt3_V214error_category10_M_messageEi .xdata$_ZNKSt3_V214error_category10_M_messageEi .pdata$_ZNKSt3_V214error_category10_M_messageEi _ZNK12_GLOBAL__N_117io_error_category4nameEv _ZN12_GLOBAL__N_122__io_category_instanceEv _ZGVZN12_GLOBAL__N_122__io_categoq	      ry_instanceEvE4__ec _ZZN12_GLOBAL__N_122__io_category_instanceEvE4__ec _ZN12_GLOBAL__N_117io_error_categoryD2Ev _ZTVN12_GLOBAL__N_117io_error_categoryE _ZN12_GLOBAL__N_117io_error_categoryD1Ev _ZN12_GLOBAL__N_117io_error_categoryD0Ev _ZNSt8ios_base7failureB5cxx11D2Ev .rdata$_ZTVNSt8ios_base7failureB5cxx11E _ZNSt8ios_base7failureB5cxx11D1Ev _ZNSt8ios_base7failureB5cxx11D0Ev _ZNKSt8ios_base7failureB5cxx114whatEv _ZNSt19__iosfail_type_infoD2Ev .rdata$_ZTVSt19__iosfail_type_info _ZNSt19__iosfail_type_infoD1Ev _ZNSt19__iosfail_type_infoD0Ev _ZNKSt19__iosfail_type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .text$_ZNSt13__ios_failureD1Ev _ZNSt13__ios_failureD1Ev .rdata$_ZTVSt13__ios_failure .text$_ZNSt13__ios_failureD0Ev _ZNSt13__ios_failureD0Ev _ZNK12_GLOBAL__N_117io_error_category7messageB5cxx11Ei _ZSt17iostream_categoryv _ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt8ios_base7failureB5cxx11C1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEEr	       _ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt10error_code _ZNSt8ios_base7failureB5cxx11C1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt10error_code _ZNSt8ios_base7failureB5cxx11C2EPKcRKSt10error_code _ZNSt8ios_base7failureB5cxx11C1EPKcRKSt10error_code _ZSt19__throw_ios_failurePKc .rdata$_ZTISt13__ios_failure .rdata$_ZTSNSt3_V214error_categoryE .rdata$_ZTINSt3_V214error_categoryE .rdata$_ZTSSt12system_error .rdata$_ZTISt12system_error .rdata$_ZTSNSt8ios_base7failureB5cxx11E .rdata$_ZTINSt8ios_base7failureB5cxx11E _ZTIN12_GLOBAL__N_117io_error_categoryE _ZTSN12_GLOBAL__N_117io_error_categoryE .rdata$_ZTSSt13__ios_failure .rdata$_ZTSSt19__iosfail_type_info .rdata$_ZTISt19__iosfail_type_info .text$_ZNK12_GLOBAL__N_117io_error_category4nameEv .xdata$_ZNK12_GLOBAL__N_117io_error_category4nameEv .pdata$_ZNK12_GLOBAL__N_117io_error_category4nameEv .text$_ZN12_GLOBAL__N_122__io_category_instanceEv .xdata$_ZN12_GLOBAL__N_122__io_category_instanceEv .pdas	      ta$_ZN12_GLOBAL__N_122__io_category_instanceEv .text$_ZN12_GLOBAL__N_117io_error_categoryD2Ev .xdata$_ZN12_GLOBAL__N_117io_error_categoryD2Ev .pdata$_ZN12_GLOBAL__N_117io_error_categoryD2Ev .text$_ZN12_GLOBAL__N_117io_error_categoryD0Ev .xdata$_ZN12_GLOBAL__N_117io_error_categoryD0Ev .pdata$_ZN12_GLOBAL__N_117io_error_categoryD0Ev .text$_ZNSt8ios_base7failureB5cxx11D2Ev .xdata$_ZNSt8ios_base7failureB5cxx11D2Ev .pdata$_ZNSt8ios_base7failureB5cxx11D2Ev .text$_ZNSt8ios_base7failureB5cxx11D0Ev .xdata$_ZNSt8ios_base7failureB5cxx11D0Ev .pdata$_ZNSt8ios_base7failureB5cxx11D0Ev .text$_ZNKSt8ios_base7failureB5cxx114whatEv .xdata$_ZNKSt8ios_base7failureB5cxx114whatEv .pdata$_ZNKSt8ios_base7failureB5cxx114whatEv .text$_ZNSt19__iosfail_type_infoD2Ev .xdata$_ZNSt19__iosfail_type_infoD2Ev .pdata$_ZNSt19__iosfail_type_infoD2Ev .text$_ZNSt19__iosfail_type_infoD0Ev .xdata$_ZNSt19__iosfail_type_infoD0Ev .pdata$_ZNSt19__iosfail_type_infoD0Ev .text$_ZNKSt19__iosfail_type_info11__do_upcastEPKN10__cxxabiv117__class_type_int	      foEPPv .xdata$_ZNKSt19__iosfail_type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .pdata$_ZNKSt19__iosfail_type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv .xdata$_ZNSt13__ios_failureD1Ev .pdata$_ZNSt13__ios_failureD1Ev .xdata$_ZNSt13__ios_failureD0Ev .pdata$_ZNSt13__ios_failureD0Ev .text$_ZNK12_GLOBAL__N_117io_error_category7messageB5cxx11Ei .xdata$_ZNK12_GLOBAL__N_117io_error_category7messageB5cxx11Ei .pdata$_ZNK12_GLOBAL__N_117io_error_category7messageB5cxx11Ei .text$_ZSt17iostream_categoryv .xdata$_ZSt17iostream_categoryv .pdata$_ZSt17iostream_categoryv .text$_ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt10error_code .xdata$_ZNSt8ios_base7failureB5cxx11Cu	      2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt10error_code .pdata$_ZNSt8ios_base7failureB5cxx11C2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEERKSt10error_code .text$_ZNSt8ios_base7failureB5cxx11C2EPKcRKSt10error_code .xdata$_ZNSt8ios_base7failureB5cxx11C2EPKcRKSt10error_code .pdata$_ZNSt8ios_base7failureB5cxx11C2EPKcRKSt10error_code .text$_ZSt19__throw_ios_failurePKc .xdata$_ZSt19__throw_ios_failurePKc .pdata$_ZSt19__throw_ios_failurePKc .rdata$_ZTIN12_GLOBAL__N_117io_error_categoryE .rdata$_ZTSN12_GLOBAL__N_117io_error_categoryE .rdata$_ZTVN12_GLOBAL__N_117io_error_categoryE .data$_ZGVZN12_GLOBAL__N_122__io_category_instanceEvE4__ec .data$_ZZN12_GLOBAL__N_122__io_category_instanceEvE4__ec _ZNSt11logic_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt11logic_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt13runtime_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt13runtime_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_trv	      aitsIcESaIcEEE _ZNSt12domain_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12domain_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt16invalid_argumentC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt16invalid_argumentC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12length_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12length_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12out_of_rangeC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12out_of_rangeC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt11range_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt11range_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt14overflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt14overflow_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt15underflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traiw	      tsIcESaIcEEE _ZNSt15underflow_errorC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12__cow_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12__cow_stringC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt11logic_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt11logic_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt11logic_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt13runtime_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt13runtime_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt13runtime_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt12domain_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt12domain_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt12domain_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt16invx	      alid_argumentC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt16invalid_argumentC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt16invalid_argumentC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt12length_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt12length_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt12length_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt12out_of_rangeC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt12out_of_rangeC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt12out_of_rangeC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt11range_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt11range_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt11range_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt14overfly	      ow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt14overflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt14overflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt15underflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt15underflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt15underflow_errorC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt12__cow_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt12__cow_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt12__cow_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12__sso_stringC2Ev _ZNSt12__sso_stringC1Ev _ZNSt12__sso_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12__sso_stringC1ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE _ZNSt12__sso_stringC2EPKcy _ZNSt12__sso_stringC1EPKcy _ZNSt12__ssz	      o_stringC2ERKS_ _ZNSt12__sso_stringC1ERKS_ _ZNSt12__sso_stringaSERKS_ _ZNSt12__sso_stringD2Ev _ZNSt12__sso_stringD1Ev _ZNSt12__sso_stringC2EOS_ _ZNSt12__sso_stringC1EOS_ _ZNSt12__sso_stringaSEOS_ .text$_ZNSt12__sso_stringC2Ev .xdata$_ZNSt12__sso_stringC2Ev .pdata$_ZNSt12__sso_stringC2Ev .text$_ZNSt12__sso_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .xdata$_ZNSt12__sso_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .pdata$_ZNSt12__sso_stringC2ERKNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEEE .text$_ZNSt12__sso_stringC2EPKcy .xdata$_ZNSt12__sso_stringC2EPKcy .pdata$_ZNSt12__sso_stringC2EPKcy .text$_ZNSt12__sso_stringC2ERKS_ .xdata$_ZNSt12__sso_stringC2ERKS_ .pdata$_ZNSt12__sso_stringC2ERKS_ .text$_ZNSt12__sso_stringaSERKS_ .xdata$_ZNSt12__sso_stringaSERKS_ .pdata$_ZNSt12__sso_stringaSERKS_ .text$_ZNSt12__sso_stringD2Ev .xdata$_ZNSt12__sso_stringD2Ev .pdata$_ZNSt12__sso_stringD2Ev .text$_ZNSt12__sso_stringC2EOS_ .xdata$_ZNSt12__sso_stringC2EOS_ .pdata$_ZNSt12__s{	      so_stringC2EOS_ .text$_ZNSt12__sso_stringaSEOS_ .xdata$_ZNSt12__sso_stringaSEOS_ .pdata$_ZNSt12__sso_stringaSEOS_ _ZNK12_GLOBAL__N_122generic_error_category4nameEv _ZNK12_GLOBAL__N_121system_error_category4nameEv _ZNKSt3_V214error_category23default_error_conditionEi _ZNKSt3_V214error_category10equivalentERKSt10error_codei _ZN12_GLOBAL__N_121system_error_categoryD2Ev _ZN12_GLOBAL__N_121system_error_categoryD1Ev _ZN12_GLOBAL__N_122generic_error_categoryD2Ev _ZN12_GLOBAL__N_122generic_error_categoryD1Ev _ZN12_GLOBAL__N_121system_error_categoryD0Ev _ZN12_GLOBAL__N_122generic_error_categoryD0Ev _ZNSt12system_errorD2Ev .rdata$_ZTVSt12system_error _ZNSt12system_errorD1Ev _ZNSt12system_errorD0Ev _ZNKSt3_V214error_category10_M_messageB5cxx11Ei _ZNK12_GLOBAL__N_122generic_error_category7messageB5cxx11Ei _ZNK12_GLOBAL__N_121system_error_category7messageB5cxx11Ei _ZNKSt3_V214error_category10equivalentEiRKSt15error_condition _ZSt20__throw_system_errori _ZN12_GLOBAL__N_1L25generic_category_instanceE _ZNSt3_V214erro|	      r_categoryD2Ev _ZNSt3_V214error_categoryD1Ev _ZNSt3_V214error_categoryD0Ev _ZNSt3_V215system_categoryEv _ZN12_GLOBAL__N_1L24system_category_instanceE _ZNSt3_V216generic_categoryEv _ZNKSt10error_code23default_error_conditionEv _GLOBAL__sub_I__ZSt20__throw_system_errori _ZTIN12_GLOBAL__N_122generic_error_categoryE _ZTSN12_GLOBAL__N_122generic_error_categoryE _ZTIN12_GLOBAL__N_121system_error_categoryE _ZTSN12_GLOBAL__N_121system_error_categoryE _ZTVN12_GLOBAL__N_122generic_error_categoryE _ZTVN12_GLOBAL__N_121system_error_categoryE .rdata$_ZTVNSt3_V214error_categoryE .text$_ZNK12_GLOBAL__N_122generic_error_category4nameEv .xdata$_ZNK12_GLOBAL__N_122generic_error_category4nameEv .pdata$_ZNK12_GLOBAL__N_122generic_error_category4nameEv .text$_ZNK12_GLOBAL__N_121system_error_category4nameEv .xdata$_ZNK12_GLOBAL__N_121system_error_category4nameEv .pdata$_ZNK12_GLOBAL__N_121system_error_category4nameEv .text$_ZNKSt3_V214error_category23default_error_conditionEi .xdata$_ZNKSt3_V214error_category23default_erro}	      r_conditionEi .pdata$_ZNKSt3_V214error_category23default_error_conditionEi .text$_ZNKSt3_V214error_category10equivalentERKSt10error_codei .xdata$_ZNKSt3_V214error_category10equivalentERKSt10error_codei .pdata$_ZNKSt3_V214error_category10equivalentERKSt10error_codei .text$_ZN12_GLOBAL__N_121system_error_categoryD2Ev .xdata$_ZN12_GLOBAL__N_121system_error_categoryD2Ev .pdata$_ZN12_GLOBAL__N_121system_error_categoryD2Ev .text$_ZN12_GLOBAL__N_122generic_error_categoryD2Ev .xdata$_ZN12_GLOBAL__N_122generic_error_categoryD2Ev .pdata$_ZN12_GLOBAL__N_122generic_error_categoryD2Ev .text$_ZN12_GLOBAL__N_121system_error_categoryD0Ev .xdata$_ZN12_GLOBAL__N_121system_error_categoryD0Ev .pdata$_ZN12_GLOBAL__N_121system_error_categoryD0Ev .text$_ZN12_GLOBAL__N_122generic_error_categoryD0Ev .xdata$_ZN12_GLOBAL__N_122generic_error_categoryD0Ev .pdata$_ZN12_GLOBAL__N_122generic_error_categoryD0Ev .text$_ZNSt12system_errorD2Ev .xdata$_ZNSt12system_errorD2Ev .pdata$_ZNSt12system_errorD2Ev .text$_ZNSt12system_errorD0Ev .x~	      data$_ZNSt12system_errorD0Ev .pdata$_ZNSt12system_errorD0Ev .text$_ZNKSt3_V214error_category10_M_messageB5cxx11Ei .xdata$_ZNKSt3_V214error_category10_M_messageB5cxx11Ei .pdata$_ZNKSt3_V214error_category10_M_messageB5cxx11Ei .text$_ZNK12_GLOBAL__N_122generic_error_category7messageB5cxx11Ei .xdata$_ZNK12_GLOBAL__N_122generic_error_category7messageB5cxx11Ei .pdata$_ZNK12_GLOBAL__N_122generic_error_category7messageB5cxx11Ei .text$__tcf_1 .xdata$__tcf_1 .pdata$__tcf_1 .text$_ZNKSt3_V214error_category10equivalentEiRKSt15error_condition .xdata$_ZNKSt3_V214error_category10equivalentEiRKSt15error_condition .pdata$_ZNKSt3_V214error_category10equivalentEiRKSt15error_condition .text$_ZSt20__throw_system_errori .xdata$_ZSt20__throw_system_errori .pdata$_ZSt20__throw_system_errori .text$_ZNSt3_V214error_categoryD2Ev .xdata$_ZNSt3_V214error_categoryD2Ev .pdata$_ZNSt3_V214error_categoryD2Ev .text$_ZNSt3_V214error_categoryD0Ev .xdata$_ZNSt3_V214error_categoryD0Ev .pdata$_ZNSt3_V214error_categoryD0Ev .text$_ZNSt3_V215s	      ystem_categoryEv .xdata$_ZNSt3_V215system_categoryEv .pdata$_ZNSt3_V215system_categoryEv .text$_ZNSt3_V216generic_categoryEv .xdata$_ZNSt3_V216generic_categoryEv .pdata$_ZNSt3_V216generic_categoryEv .text$_ZNKSt10error_code23default_error_conditionEv .xdata$_ZNKSt10error_code23default_error_conditionEv .pdata$_ZNKSt10error_code23default_error_conditionEv .text.startup._GLOBAL__sub_I__ZSt20__throw_system_errori .xdata.startup._GLOBAL__sub_I__ZSt20__throw_system_errori .pdata.startup._GLOBAL__sub_I__ZSt20__throw_system_errori .rdata$_ZTIN12_GLOBAL__N_122generic_error_categoryE .rdata$_ZTSN12_GLOBAL__N_122generic_error_categoryE .rdata$_ZTIN12_GLOBAL__N_121system_error_categoryE .rdata$_ZTSN12_GLOBAL__N_121system_error_categoryE .rdata$_ZTVN12_GLOBAL__N_122generic_error_categoryE .rdata$_ZTVN12_GLOBAL__N_121system_error_categoryE .data$_ZN12_GLOBAL__N_1L24system_category_instanceE .data$_ZN12_GLOBAL__N_1L25generic_category_instanceE _ZNSi6ignoreEx _ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEx .text$�	      _ZNSi6ignoreEx .xdata$_ZNSi6ignoreEx .pdata$_ZNSi6ignoreEx .text$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEx .xdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEx .pdata$_ZNSt13basic_istreamIwSt11char_traitsIwEE6ignoreEx _ZNKSt20bad_array_new_length4whatEv _ZNSt20bad_array_new_lengthD2Ev .rdata$_ZTVSt20bad_array_new_length _ZNSt20bad_array_new_lengthD1Ev _ZNSt20bad_array_new_lengthD0Ev .text$_ZNKSt20bad_array_new_length4whatEv .xdata$_ZNKSt20bad_array_new_length4whatEv .pdata$_ZNKSt20bad_array_new_length4whatEv .text$_ZNSt20bad_array_new_lengthD2Ev .xdata$_ZNSt20bad_array_new_lengthD2Ev .pdata$_ZNSt20bad_array_new_lengthD2Ev .text$_ZNSt20bad_array_new_lengthD0Ev .xdata$_ZNSt20bad_array_new_lengthD0Ev .pdata$_ZNSt20bad_array_new_lengthD0Ev d_make_comp d_ref_qualifier d_count_templates_scopes d_append_buffer d_number.isra.0 d_number_component d_compact_number d_template_param d_source_name d_abi_tags d_substitution standard_subs d_call_offset next_is_type_qual.isra.2 d_discriminator d_index_t�	      emplate_argument.part.8 d_lookup_template_argument.isra.9 d_find_pack d_growable_string_callback_adapter d_expr_primary d_expression_1 d_exprlist d_template_args_1 d_template_args cplus_demangle_builtin_types d_type.cold.23 d_operator_name cplus_demangle_operators d_parmlist d_cv_qualifiers d_bare_function_type d_function_type d_unqualified_name CSWTCH.125 d_encoding d_print_comp_inner d_print_comp d_print_mod d_print_function_type.isra.14 d_print_mod_list d_print_array_type.isra.13 d_print_expr_op d_print_subexpr d_maybe_print_fold_expression.isra.19 d_demangle_callback.constprop.21 __cxa_demangle __gcclibcxx_demangle_callback .text.unlikely .xdata.unlikely .pdata.unlikely __cxa_call_terminate .text$__cxa_call_terminate .xdata$__cxa_call_terminate .pdata$__cxa_call_terminate __cxa_current_exception_type .text$__cxa_current_exception_type .xdata$__cxa_current_exception_type .pdata$__cxa_current_exception_type _ZnwyRKSt9nothrow_t .text$_ZnwyRKSt9nothrow_t .xdata$_ZnwyRKSt9nothrow_t .pdata$_ZnwyRKSt9not�	      hrow_t _ZNKSt8ios_base7failure4whatEv _ZNSt8ios_base7failureD2Ev .rdata$_ZTVNSt8ios_base7failureE _ZNSt8ios_base7failureD1Ev _ZNSt8ios_base7failureD0Ev _ZNSt8ios_base7failureC2ERKSs _ZNSt8ios_base7failureC1ERKSs _ZSt23__construct_ios_failurePvPKc _ZSt21__destroy_ios_failurePv _ZSt24__is_ios_failure_handlerPKN10__cxxabiv117__class_type_infoE .rdata$_ZTINSt8ios_base7failureE .rdata$_ZTSNSt8ios_base7failureE .text$_ZNKSt8ios_base7failure4whatEv .xdata$_ZNKSt8ios_base7failure4whatEv .pdata$_ZNKSt8ios_base7failure4whatEv .text$_ZNSt8ios_base7failureD2Ev .xdata$_ZNSt8ios_base7failureD2Ev .pdata$_ZNSt8ios_base7failureD2Ev .text$_ZNSt8ios_base7failureD0Ev .xdata$_ZNSt8ios_base7failureD0Ev .pdata$_ZNSt8ios_base7failureD0Ev .text$_ZNSt8ios_base7failureC2ERKSs .xdata$_ZNSt8ios_base7failureC2ERKSs .pdata$_ZNSt8ios_base7failureC2ERKSs .text$_ZSt23__construct_ios_failurePvPKc .xdata$_ZSt23__construct_ios_failurePvPKc .pdata$_ZSt23__construct_ios_failurePvPKc .text$_ZSt21__destroy_ios_failurePv .xdata$_ZSt21__destro�	      y_ios_failurePv .pdata$_ZSt21__destroy_ios_failurePv .text$_ZSt24__is_ios_failure_handlerPKN10__cxxabiv117__class_type_infoE .xdata$_ZSt24__is_ios_failure_handlerPKN10__cxxabiv117__class_type_infoE .pdata$_ZSt24__is_ios_failure_handlerPKN10__cxxabiv117__class_type_infoE __do_global_dtors __do_global_ctors .rdata$.refptr.__CTOR_LIST__ initialized my_lconv_init __security_init_cookie .data$__security_cookie .data$__security_cookie_complement __report_gsfailure GS_ContextRecord GS_ExceptionRecord GS_ExceptionPointers __dyn_tls_dtor __dyn_tls_init .rdata$.refptr._CRT_MT __tlregdtor __mingw_raise_matherr stUserMathErr __mingw_setusermatherr _decode_pointer _encode_pointer __report_error __write_memory.part.0 maxSections _pei386_runtime_relocator was_init.95174 .rdata$.refptr.__RUNTIME_PSEUDO_RELOC_LIST_END__ .rdata$.refptr.__RUNTIME_PSEUDO_RELOC_LIST__ __mingw_SEH_error_handler __mingw_init_ehandler was_here.95013 emu_pdata emu_xdata _gnu_exception_handler __mingwthr_run_key_dtors.part.0 __mingwthr_cs key_�	      dtor_list ___w64_mingwthr_add_key_dtor __mingwthr_cs_init ___w64_mingwthr_remove_key_dtor __mingw_TLScallback pseudo-reloc-list.c _ValidateImageBase.part.0 _ValidateImageBase _FindPESection _FindPESectionByName __mingw_GetSectionForAddress __mingw_GetSectionCount _FindPESectionExec _GetPEImageBase _IsNonwritableInCurrentImage __mingw_enum_import_library_names _Unwind_ForcedUnwind_Phase2 _Unwind_GetGR _Unwind_SetGR _Unwind_GetCFA _Unwind_GetIP _Unwind_GetIPInfo _Unwind_SetIP _Unwind_GetLanguageSpecificData _Unwind_GetRegionStart _Unwind_FindEnclosingFunction _Unwind_GetDataRelBase _Unwind_GetTextRelBase _GCC_specific_handler _Unwind_RaiseException _Unwind_Resume _Unwind_Resume_or_Rethrow _Unwind_ForcedUnwind _Unwind_DeleteException _Unwind_Backtrace .debug_loc emutls_destroy emutls_init emutls_mutex emutls_key __emutls_get_address once.8585 emutls_size __emutls_register_common .debug_ranges __mingw_strtod fpi0.4260 __mingw_strtof __mbrtowc_cp internal_mbstate.53756 mbsrtowcs internal_mbstate.53767 s_mb�	      state.53783 __asctoe64 __wcrtomb_cp wcsrtombs _ftelli64 .rdata$.refptr.__imp___pioinfo _fseeki64 mingw_dosmaperr local_errtab __mingw_vsnprintf __increment_D2A __decrement_D2A __set_ones_D2A __strtodg .rdata$.refptr.__tens_D2A fivesbits .rdata$.refptr.__bigtens_D2A .rdata$.refptr.__tinytens_D2A __sum_D2A __eshift.part.3 __enormlz __emdnorm __pformat_cvt __pformat_putc __pformat_wputchars __pformat_putchars __pformat_puts __pformat_emit_inf_or_nan __pformat_emit_radix_point __pformat_emit_float __pformat_float __pformat_int.isra.0 __pformat_emit_efloat __pformat_efloat __pformat_gfloat __pformat_xint.isra.1 __pformat_xldouble __mingw_pformat __rv_alloc_D2A __nrv_alloc_D2A __freedtoa __quorem_D2A __gethex_D2A .rdata$.refptr.__hexdig_D2A __rshift_D2A __trailz_D2A __mingw_hexdig_init_D2A __hexnan_D2A dtoa_lock dtoa_CS_init dtoa_CritSec dtoa_lock_cleanup __Balloc_D2A pmem_next private_mem __Bfree_D2A __multadd_D2A __i2b_D2A __mult_D2A __pow5mult_D2A p05.53702 __lshift_D2A __cmp_D2A __diff_D2A __b2d_D2A __d�	      2b_D2A __strcp_D2A __s2b_D2A __ratio_D2A __match_D2A __copybits_D2A __any_on_D2A __acrt_iob_func mingw_get_invalid_parameter_handler _get_invalid_parameter_handler mingw_set_invalid_parameter_handler _set_invalid_parameter_handler invalid_parameter_handler.c __p__acmdln .rdata$.refptr.__imp__acmdln __p__fmode .rdata$.refptr.__imp__fmode do_sema_b_release cond_print_set print_state cond_print pthread_condattr_destroy pthread_condattr_init pthread_condattr_getpshared pthread_condattr_getclock pthread_condattr_setclock __pthread_clock_nanosleep pthread_condattr_setpshared pthread_cond_init cond_static_init cond_locked do_sema_b_wait_intern do_sema_b_wait pthread_cond_destroy pthread_cond_signal pthread_cond_broadcast pthread_cond_wait cleanup_wait pthread_cond_timedwait_impl pthread_cond_timedwait pthread_cond_timedwait_relative_np _pthread_time_in_ms _pthread_time_in_ms_from_timespec _pthread_rel_time_in_ms mutex_impl_init pthread_mutex_lock pthread_mutex_timedlock pthread_mutex_unlock pthread_mutex_try�	      lock pthread_mutex_init pthread_mutex_destroy pthread_mutexattr_init pthread_mutexattr_destroy pthread_mutexattr_gettype pthread_mutexattr_settype pthread_mutexattr_getpshared pthread_mutexattr_setpshared pthread_mutexattr_getprotocol pthread_mutexattr_setprotocol pthread_mutexattr_getprioceiling pthread_mutexattr_setprioceiling pthread_spin_init pthread_spin_destroy pthread_spin_lock pthread_spin_trylock pthread_spin_unlock SetThreadName_VEH enterOnceObject once_global pthread_tls_init _pthread_tls __pthread_get_pointer idListCnt __pthread_register_pointer idListMax idListNextId push_pthread_mem.part.2 mtx_pthr_locked pthr_last pthr_root leaveOnceObject.part.4 _pthread_once_cleanup pop_pthread_mem replace_spin_keys.constprop.10 _pthread_once_raw.part.5.constprop.11 _pthread_tls_once __pthread_self_lite __pth_gpointer_locked _pthread_cleanup_dest.part.8 _pthread_key_lock __dyn_tls_pthread SetThreadName_VEH_handle pthread_create_wrapper .tl_start thread_print_set thread_print pthread_timechange_handler�	      _np pthread_num_processors_np pthread_set_num_processors_np pthread_once pthread_key_create _pthread_key_sch _pthread_key_max pthread_key_delete pthread_getspecific pthread_setspecific pthread_equal _pthread_cleanup_dest pthread_self pthread_getevent pthread_gethandle pthread_getclean pthread_get_concurrency _pthread_concur pthread_set_concurrency pthread_exit __pthread_shallcancel _pthread_cancelling _pthread_setnobreak _pthread_invoke_cancel test_cancel_locked pthread_testcancel pthread_delay_np pthread_delay_np_ms pthread_cancel pthread_kill _pthread_get_state _pthread_set_state pthread_attr_init pthread_attr_destroy pthread_attr_setdetachstate pthread_attr_getdetachstate pthread_attr_setinheritsched pthread_attr_getinheritsched pthread_attr_setscope pthread_attr_getscope pthread_attr_getstackaddr pthread_attr_setstackaddr pthread_attr_getstacksize pthread_attr_setstacksize pthread_setcancelstate pthread_setcanceltype pthread_create pthread_join _pthread_tryjoin pthread_detach pthread_getconcurrenc�	      y dummy_concurrency_level pthread_setconcurrency pthread_setname_np pthread_getname_np rwl_ref_destroy rwl_global rwl_ref_unlock rwlock_gain_both_locks rwlock_free_both_locks st_cancelwrite rwl_unref rwl_print_set rwl_print pthread_rwlock_init rwlock_static_init rwl_ref.isra.0 pthread_rwlock_destroy pthread_rwlock_rdlock pthread_rwlock_timedrdlock pthread_rwlock_tryrdlock pthread_rwlock_trywrlock pthread_rwlock_unlock pthread_rwlock_wrlock pthread_rwlock_timedwrlock pthread_rwlockattr_destroy pthread_rwlockattr_init pthread_rwlockattr_getpshared pthread_rwlockattr_setpshared mingw_getsp register_frame_ctor .text.startup .xdata.startup .pdata.startup .ctors.65535 _ZTSN10__cxxabiv115__forced_unwindE _ZTSSt14basic_iostreamIwSt11char_traitsIwEE __imp___acrt_iob_func _ZTVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .refptr._ZTVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZTISt13basic_filebufIcSt11char_traitsIcEE .refptr._ZTVSt15underflow_error _ZTVN10__cxxab�	      iv120__si_class_type_infoE _ZTVSt15numpunct_bynameIwE _ZN14__gnu_internal7buf_cinE .refptr._ZNSt10moneypunctIwLb0EE2idE __imp_CreateSemaphoreA _dowildcard _ZTSSt8messagesIcE _ZTIN10__cxxabiv115__forced_unwindE _ZTINSt7__cxx1110moneypunctIcLb0EEE __imp_Sleep _ZTISt18__moneypunct_cacheIwLb1EE __imp_EnterCriticalSection _ZTSSt13basic_filebufIcSt11char_traitsIcEE _ZTSSt21__ctype_abstract_baseIwE _ZNSt8ios_base6binaryE .refptr.__hexdig_D2A .refptr.__RUNTIME_PSEUDO_RELOC_LIST__ __imp_memcmp .refptr._ZTVSt11range_error _ZTISt13bad_exception _ZTVSt12length_error _ZNSt10ctype_base5digitE _ZTVSt12system_error _ZTINSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE __imp_strcoll _ZTVSt15messages_bynameIwE _ZTISt7codecvtIwciE CloseHandle .refptr._ZTVSt12domain_error __imp_read _ZTVSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTSSt15basic_streambufIwSt11char_traitsIwEE _ZTISt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZTSSt7collateIwE .refptr._ZN10__cxxabiv119__termin�	      ate_handlerE _ZTISt18__moneypunct_cacheIcLb1EE _ZTVSt10moneypunctIcLb0EE GetCurrentProcess __imp__endthreadex SetProcessAffinityMask GetCurrentProcessId __imp_strlen _ZNSt17moneypunct_bynameIcLb1EE4intlE __imp_malloc __imp___getmainargs ___crt_xi_end__ _ZTVN10__cxxabiv117__class_type_infoE _ZN14__gnu_internal8buf_cerrE _ZTISt21__ctype_abstract_baseIcE _ZTTSt13basic_ostreamIwSt11char_traitsIwEE mingw_pcinit _ZTISt16invalid_argument __imp_VirtualQuery __imp__fmode _ZTVNSt7__cxx1117moneypunct_bynameIwLb1EEE _ZTCSt14basic_ofstreamIcSt11char_traitsIcEE0_So .refptr._gnu_exception_handler _ZNSt10ctype_base5upperE .refptr._ZNSt10bad_typeidD1Ev .refptr._ZNSt7__cxx118numpunctIcE2idE _ZNSt6locale5_Impl11_S_id_ctypeE _ZNSt10ctype_base5spaceE _ZNSt7__cxx118messagesIcE2idE .refptr._ZSt4cerr _ZTISt19__codecvt_utf8_baseIwE .refptr._ZTVNSt7__cxx117collateIcEE __tens_D2A .refptr._ZNSt7__cxx117collateIwE2idE GetThreadContext .refptr._ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp_GetHandleInforma�	      tion _ZNSt6locale4timeE __imp_RtlAddFunctionTable _ZTVSt16__numpunct_cacheIwE __rt_psrelocs_start __imp__filelengthi64 _strnicmp .refptr._ZNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE __IAT_end__ .refptr._matherr _ZTISt17moneypunct_bynameIcLb1EE _ZNSt8ios_base10scientificE AddVectoredExceptionHandler __imp_sprintf _ZNSt8ios_base4Init20_S_synced_with_stdioE _ZTIN9__gnu_cxx24__concurrence_lock_errorE _ZTSNSt7__cxx1114collate_bynameIwEE __imp_fprintf _ZTVSt12domain_error _ZNSt8messagesIwE2idE _ZTSNSt7__cxx118messagesIcEE _ZTSSt19__iosfail_type_info _ZGVNSt7collateIcE2idE _ZGVNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr._ZNSt12length_errorD1Ev .refptr._CRT_MT _ZTINSt7__cxx1114collate_bynameIcEE _ZGVNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt5ctypeIwE _ZTVSt18__moneypunct_cacheIcLb1EE _ZTVNSt7__cxx117collateIwEE .refptr._ZSt5wcerr _ZNSt7__cxx119money_p�	      utIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE SuspendThread CreateSemaphoreA _ZTIN10__cxxabiv119__foreign_exceptionE _ZTSSt23__codecvt_abstract_baseIcciE _ZGVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZNSt7__cxx1110moneypunctIwLb1EE2idE ___RUNTIME_PSEUDO_RELOC_LIST_END__ _ZNSt8ios_base11adjustfieldE _ZTISt12length_error __imp_SuspendThread _ZGVNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt8numpunctIwE2idE _ZNSt8ios_base9uppercaseE _ZTINSt8ios_base7failureE __imp_CloseHandle _ZTISt9exception .refptr._ZTVSt7collateIwE _ZNSt7collateIcE2idE _ZTISt13basic_fstreamIwSt11char_traitsIwEE _ZTISt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE RemoveVectoredExceptionHandler _ZNSt10__num_base12_S_atoms_outE _ZTISt11logic_error _ZTVSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt15numpunct_bynameIcE _ZN14__gnu_internal13buf_cerr_syncE .refptr._ZSt3cin .refptr._ZN14__gnu_internal9buf_wcoutE _ZTINSt7__cxx1110moneypunctIwLb0E�	      EE __imp_SetLastError SetThreadPriority ___crt_xc_start__ __imp___setusermatherr _ZTISt7codecvtIDiciE _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE __imp_strxfrm _ZTISt15numpunct_bynameIcE __imp_strdup .refptr._ZTVSt14overflow_error _ZTCSt13basic_fstreamIwSt11char_traitsIwEE0_St13basic_istreamIwS1_E .refptr._ZNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr.__imp___initenv _ZTSSt20bad_array_new_length _ZTSN10__cxxabiv117__class_type_infoE .refptr._ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr.__CTOR_LIST__ _ZTVSt7collateIwE _ZTVSt8ios_base _ZTVSt18__moneypunct_cacheIwLb1EE .refptr._ZTVSt17__timepunct_cacheIcE _ZTSSt10moneypunctIwLb0EE _ZNSt6locale5_Impl10_S_id_timeE _ZTSSt25__codecvt_utf8_utf16_baseIDsE _ZTVSt11range_error _ZTSSt8ios_base _ZTSSt11range_error __imp_DuplicateHandle __hexdig_D2A _ZTSN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE _ZNSt8ios_base6eofbitE .refptr._ZNSt8ios_base4Init11_S_refcountE _ZTVSt14basi�	      c_ifstreamIwSt11char_traitsIwEE _ZGVNSt10moneypunctIcLb0EE2idE .refptr._ZTVSt18__moneypunct_cacheIcLb0EE .refptr._ZN14__gnu_internal8buf_cerrE _ZTVSt7codecvtIDiciE __imp_DeleteCriticalSection __imp_OutputDebugStringA __major_os_version__ _ZNSt8ios_base4leftE _ZTVSt18__moneypunct_cacheIwLb0EE _ZTVSt20__codecvt_utf16_baseIwE .refptr._ZTVSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt14codecvt_bynameIcciE _ZTVSt7collateIcE __imp__set_invalid_parameter_handler _ZTINSt7__cxx1115numpunct_bynameIcEE _ZTSSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt5ctypeIcE .refptr.__image_base__ _ZTSSt9basic_iosIwSt11char_traitsIwEE _ZTSNSt7__cxx1117moneypunct_bynameIcLb1EEE .refptr._ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt12domain_error _ZTSN10__cxxabiv120__si_class_type_infoE __imp_GetThreadPriority _ZTSN9__gnu_cxx26__concurrence_unlock_errorE _ZTSNSt7__cxx118numpunctIcEE _ZTVSt13basic_filebufIwSt11char_traitsIwEE _ZTVSt17moneypunct_bynameIcLb0EE __imp_f�	      puts _ZTVNSt7__cxx1117moneypunct_bynameIwLb0EEE _ZTSSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTIN9__gnu_cxx29__concurrence_broadcast_errorE __doserrno _ZTSSt12codecvt_base _ZTSSt19__codecvt_utf8_baseIDiE _ZTSSt13bad_exception __imp_calloc __imp__fileno .refptr._ZSt4clog .refptr._ZTVSt16invalid_argument _ZTTSt14basic_ofstreamIwSt11char_traitsIwEE __imp_GetThreadContext _ZGVNSt7__cxx118numpunctIwE2idE .refptr._ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE __loader_flags__ .refptr._newmode __size_of_heap_commit__ _ZTISt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt17moneypunct_bynameIwLb0EE4intlE _ZNSt7__cxx117collateIwE2idE _ZNSt7codecvtIDsciE2idE __C_specific_handler _ZNSt8ios_base5truncE .refptr.mingw_initcharmax _ZTSSt18__moneypunct_cacheIwLb0EE .refptr._ZNSt13bad_exceptionD1Ev _ZNSt10money_base18_S_default_patternE _ZTSNSt7__cxx1114collate_bynameIcEE __imp_RtlVirtualUnwind .refptr._ZTVSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _�	      _imp_GetTickCount __imp_strftime _ZTISt12ctype_bynameIcE _ZTISt19__codecvt_utf8_baseIDsE __RUNTIME_PSEUDO_RELOC_LIST__ __imp__amsg_exit _ZNSt8ios_base7failbitE _ZTISt8numpunctIwE .refptr._ZTVNSt7__cxx1110moneypunctIcLb0EEE __imp_memcpy _ZTISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE __imp__strnicmp _ZNSt8ios_base9showpointE _ZTISt8messagesIcE _ZTVSt8messagesIwE _ZTSSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZTISt20__codecvt_utf16_baseIwE ResetEvent _ZTCSt14basic_iostreamIwSt11char_traitsIwEE16_St13basic_ostreamIwS1_E .refptr._ZTVSt10moneypunctIcLb0EE .refptr._ZTVSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt13basic_fstreamIwSt11char_traitsIwEE __imp_fdopen _ZTSSt17moneypunct_bynameIcLb1EE __mingw_winmain_nShowCmd _ZTISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt9basic_iosIcSt11char_traitsIcEE _ZNSt7__cxx1110moneypunctIwLb1EE2idE IsDebuggerPresent __imp_strtoul _ZTSSt18__moneypunct_cacheIcLb1EE .refptr._ZNSt5ctypeIwE2idE .refptr�	      ._ZN14__gnu_internal13buf_cerr_syncE _ZTISt8messagesIwE _ZTSSt16__numpunct_cacheIwE __rt_psrelocs_size _ZTSSt16invalid_argument _ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt10moneypunctIwLb1EE .refptr._ZTVSt17__timepunct_cacheIwE TerminateProcess .refptr._ZNSt10money_base8_S_atomsE _ZTISt13basic_filebufIwSt11char_traitsIwEE _ZNSt5ctypeIwE2idE __security_cookie _ZTVSt19__iosfail_type_info .refptr._ZNSt6locale9_S_globalE _ZGVNSt7__cxx117collateIwE2idE _ZNSt6locale5ctypeE _ZTINSt3_V214error_categoryE __imp_SetThreadContext __imp__get_invalid_parameter_handler .refptr._ZTVSt7codecvtIDiciE _ZNSt6locale5_Impl14_S_id_monetaryE .refptr._ZNSt7__cxx1110moneypunctIcLb1EE2idE __imp_TlsGetValue ReleaseSemaphore .refptr._ZTVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .refptr._ZTVSt14codecvt_bynameIwciE _ZTSSt17moneypunct_bynameIwLb1EE .refptr._ZNSt12domain_errorD1Ev .refptr.__imp__fmode _ZTVSt15basic_streambufIcSt11char_traitsIcEE _ZTSNSt7__cxx117collate�	      IwEE IsDBCSLeadByteEx GetCurrentThread _ZTISt13basic_ostreamIwSt11char_traitsIwEE _ZNSt8numpunctIcE2idE __imp_fileno _ZTSSt14basic_ofstreamIcSt11char_traitsIcEE _ZTIN10__cxxabiv117__class_type_infoE _ZNSt7__cxx1117moneypunct_bynameIwLb1EE4intlE _ZGVNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt10moneypunctIcLb0EE2idE _ZNSt10ctype_base5alnumE _ZN14__gnu_internal9buf_wcoutE TlsGetValue _amsg_exit _ZTVSt12out_of_range _ZTIN9__gnu_cxx24__concurrence_wait_errorE _ZTVNSt7__cxx118numpunctIwEE _ZNSt10ctype_base5printE _ZN10__cxxabiv120__unexpected_handlerE mingw_app_type _ZNSt6locale13_S_categoriesE _ZTISt7collateIwE _ZNSt7__cxx1112basic_stringIcSt11char_traitsIcESaIcEE4nposE __native_dllmain_reason __set_app_type _ZNSt8ios_base3begE _ZTVN9__gnu_cxx26__concurrence_unlock_errorE _ZTISt13__ios_failure .refptr._ZN14__gnu_internal9buf_wcerrE _ZTINSt7__cxx1114collate_bynameIwEE _ZGVNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp__lseeki64 .refptr._ZTVSt12out_of_range _ZTI�	      N10__cxxabiv120__si_class_type_infoE _ZTSNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE _ZTVNSt7__cxx1110moneypunctIwLb1EEE _ZTISt10moneypunctIcLb0EE __imp_SetUnhandledExceptionFilter mingw_pcppinit .refptr._ZTVSt7collateIcE WideCharToMultiByte __imp_RtlLookupFunctionEntry _ZTVNSt6locale5facetE _ZNSt7__cxx1110moneypunctIcLb0EE4intlE .refptr._ZSt4wcin _ZTSSt9type_info __imp_memchr _ZTSSt20__codecvt_utf16_baseIDiE _ZTVSt11logic_error _ZTVSt9exception __imp__acmdln _ZTSSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZNSt8numpunctIwE2idE _ZNSt8ios_base3outE __imp__beginthreadex _ZNSt7__cxx1110moneypunctIcLb1EE2idE _ZTVSt17moneypunct_bynameIwLb1EE _ZTIN9__gnu_cxx26__concurrence_unlock_errorE _ZTVNSt7__cxx1115numpunct_bynameIcEE .refptr._ZN14__gnu_internal13buf_wcin_syncE .refptr._ZTVNSt7__cxx118numpunctIwEE _ZTSSt12out_of_range .refptr._ZTVSt10moneypunctIwLb1EE _ZNSt8time_putIcSt19ostreambuf_iteratorI�	      cSt11char_traitsIcEEE2idE __imp_RemoveVectoredExceptionHandler __tinytens_D2A .refptr.__xc_a _ZTVSt9basic_iosIcSt11char_traitsIcEE _ZTSSt20__codecvt_utf16_baseIwE _ZTVSt14codecvt_bynameIwciE _ZTVNSt7__cxx1117moneypunct_bynameIcLb0EEE QueryPerformanceCounter _ZTTSt13basic_istreamIwSt11char_traitsIwEE _ZGVNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp_QueryPerformanceCounter _ZTSSt13basic_fstreamIcSt11char_traitsIcEE _ZGVNSt10moneypunctIcLb1EE2idE _ZNSt17__timepunct_cacheIcE12_S_timezonesE .refptr._ZTVNSt7__cxx118numpunctIcEE _ZTSNSt7__cxx1110moneypunctIwLb0EEE __imp_iswctype __imp_IsDebuggerPresent .refptr._ZNSt10money_base18_S_default_patternE _ZTSSt13messages_base _ZTVSt15basic_streambufIwSt11char_traitsIwEE _ZTVSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZSt4cerr .refptr._MINGW_INSTALL_DEBUG_MATHERR _ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp_wcslen _ZTVN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE _ZNSt10moneypu�	      nctIwLb0EE2idE _ZTSSt14codecvt_bynameIcciE _ZTVN9__gnu_cxx24__concurrence_lock_errorE .refptr.mingw_initltssuo_force _ZTINSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE EnterCriticalSection _ZN14__gnu_internal13buf_wcin_syncE _ZTSNSt7__cxx1110moneypunctIcLb1EEE .refptr.__tens_D2A _ZN14__gnu_internal8buf_coutE _ZTSSt7codecvtIDsciE _ZTSSt9bad_alloc _ZTINSt7__cxx1110moneypunctIwLb1EEE _ZGVNSt7__cxx1110moneypunctIwLb1EE2idE .refptr._ZTVSt12length_error .refptr._ZN14__gnu_internal14buf_wcout_syncE _ZNSt7codecvtIcciE2idE _tls_used _ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Si _ZGVNSt7__cxx1110moneypunctIwLb0EE2idE _ZTVSt8numpunctIcE .refptr.__bigtens_D2A _ZTISt14basic_ofstreamIwSt11char_traitsIwEE _ZTISt20__codecvt_utf16_baseIDiE GetStartupInfoA _ZTVNSt7__cxx117collateIcEE .refptr._ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE __native_startup_lock __RUNTIME_PSEUDO_RELOC_LIST_END__ _ZNSt6locale5_Impl13_S_id_numericE _ZTSSt5ctypeIcE _ZN14__gnu_internal14buf_wcout_sy�	      ncE _ZTTSt14basic_iostreamIwSt11char_traitsIwEE .refptr._ZTVSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZTSSt13basic_fstreamIwSt11char_traitsIwEE ___tls_end__ _beginthreadex .refptr._ZNSt17__timepunct_cacheIcE12_S_timezonesE __image_base__ _ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTVSt20__codecvt_utf16_baseIDsE .refptr._ZNSt17__timepunct_cacheIwE12_S_timezonesE ___crt_xp_start__ _ZTVSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE __imp_wcscoll WaitForSingleObject _ZTSSt13__ios_failure _ZTVSt25__codecvt_utf8_utf16_baseIwE _ZTVSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE OutputDebugStringA .refptr._ZTVN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE _ZTVSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE __imp_GetCurrentThreadId .refptr.__xc_z _ZGVNSt8numpunctIwE2idE _ZNSt6locale5facet7_S_onceE __imp_GetStartupInfoA _ZTVSt8bad_cast __imp_longjmp _ZTSSt10bad_typeid _ZSt4wcin _ZTSSt15numpunct_bynameIwE _ZTVSt7c�	      odecvtIwciE _ZTVSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr._ZTVSt23__codecvt_abstract_baseIcciE __imp_GetProcessAffinityMask _ZGVNSt7__cxx1110moneypunctIcLb1EE2idE _ZTISt14overflow_error .refptr._ZNSt6locale10_S_classicE __imp___lconv_init _ZTSSt11__timepunctIcE __imp_WaitForSingleObject .refptr._ZNSt7__cxx1110moneypunctIcLb0EE2idE _ZTVSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE __imp_TlsAlloc __imp_SetThreadPriority _ZN10__cxxabiv119__terminate_handlerE _ZTSSt8messagesIwE _ZTSSt10moneypunctIcLb0EE _ZNSt6locale3allE .refptr._ZNSt7__cxx1110moneypunctIwLb0EE2idE SetThreadContext _ZNSt10ctype_base5graphE __imp_fread __imp_write _ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Sd _ZTSSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZTVSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .refptr._ZNSt7__cxx118messagesIcE2idE .refptr._ZNSt7codecvtIDsciE2idE .re�	      fptr._ZTVSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE __imp_abort _ZTSSt14basic_ifstreamIwSt11char_traitsIwEE _ZTSN10__cxxabiv121__vmi_class_type_infoE _ZTSSt11__timepunctIwE _ZNSs4nposE _ZTVSt25__codecvt_utf8_utf16_baseIDiE __imp_towlower .refptr._ZNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZTVSt21__ctype_abstract_baseIwE __imp__cexit _ZTISt7collateIcE __imp_WideCharToMultiByte SetUnhandledExceptionFilter _ZTVSt19__codecvt_utf8_baseIwE _ZTINSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE ___DTOR_LIST__ .refptr._ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .refptr._ZNSt7collateIcE2idE _ZTSNSt7__cxx117collateIcEE .refptr._ZNSt7__cxx118numpunctIwE2idE _ZNSt7__cxx117collateIcE2idE _ZSt4cout __native_startup_state _head_lib64_libmsvcrt_os_a _ZTVSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTSSt12domain_error _ZTINSt�	      7__cxx1117moneypunct_bynameIcLb1EEE _ZTISt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZN14__gnu_internal9buf_wcerrE _ZSt7nothrow _ZNSt8ios_base8internalE .refptr._fmode _ZTSSt13basic_ostreamIwSt11char_traitsIwEE _ZTINSt7__cxx1115messages_bynameIwEE .refptr._ZTVSt13basic_ostreamIwSt11char_traitsIwEE __imp_wcsxfrm _ZTSSt12length_error _ZTVN9__gnu_cxx29__concurrence_broadcast_errorE __rt_psrelocs_end _ZTCSd16_So GetThreadPriority __imp_SetProcessAffinityMask __imp_getwc _ZNSt8ios_base3ateE _ZTVSt14basic_ifstreamIcSt11char_traitsIcEE _ZTTSt13basic_fstreamIwSt11char_traitsIwEE _ZTVNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE _ZTISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVN9__gnu_cxx24__concurrence_wait_errorE _ZTINSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE _ZTVNSt8ios_base7failureE _ZTISt12system_error _ZGVNSt11__timepunctIwE2idE ResumeThread __iob_func _�	      ZTVSt16invalid_argument _ZTVSt10moneypunctIcLb1EE _ZNSt11__timepunctIwE2idE _ZTSSt5ctypeIwE _ZN14__gnu_internal14buf_wcerr_syncE _ZNSt7__cxx1112basic_stringIwSt11char_traitsIwESaIwEE4nposE _ZTISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTSSt15numpunct_bynameIcE _ZTVNSt7__cxx1110moneypunctIcLb0EEE __imp_free _ZTISt10bad_typeid __imp_RaiseException _ZTISt15basic_streambufIwSt11char_traitsIwEE __imp_setlocale RtlVirtualUnwind .refptr._ZTVSt8numpunctIcE _ZNSt8ios_base6badbitE _ZTVN10__cxxabiv119__foreign_exceptionE _ZTSSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZTVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .refptr._ZTVSt13runtime_error _ZTVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _endthreadex __imp_GetCurrentThread _ZTISt25__codecvt_utf8_utf16_baseIwE __imp_WaitForMultipleObjects .refptr._ZNSt10__num_base12_S_atoms_outE ___mb_cur_max_func _ZTSSt7collateIcE _ZTINSt7__cxx118messagesIcEE .refptr._ZNSt9money_putIw�	      St19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTIN10__cxxabiv121__vmi_class_type_infoE _ZTVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZTSSt18__moneypunct_cacheIwLb1EE .refptr._ZNSt8numpunctIcE2idE _ZTISt18__moneypunct_cacheIcLb0EE _ZTINSt6locale5facet6__shimE _ZTINSt7__cxx117collateIcEE __security_cookie_complement _ZTVSt7codecvtIcciE _ZTSSt7codecvtIcciE _ZTSSt9exception _ZTINSt7__cxx1110moneypunctIcLb1EEE _ZTVSt13basic_fstreamIcSt11char_traitsIcEE _ZNSs4_Rep11_S_max_sizeE __imp_TryEnterCriticalSection _ZTVN10__cxxabiv121__vmi_class_type_infoE _ZTVSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZTVSt13runtime_error __imp_LeaveCriticalSection _ZTSSt12system_error _ZNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt25__codecvt_utf8_utf16_baseIDiE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE __imp___set_app_type _ZTISt10ctype_base __minor_subsystem_version__ _ZTVNSt7__cxx118messagesIcEE _ZNSt6locale5_Impl13_S_id_colla�	      teE _ZNSt10money_base8_S_atomsE __size_of_heap_reserve__ _ZTINSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE .refptr._ZTVSt7codecvtIDsciE .refptr._ZTVSt9basic_iosIwSt11char_traitsIwEE _ZGVNSt7__cxx117collateIcE2idE _ZTVSt19__codecvt_utf8_baseIDsE _ZTVSt13bad_exception _ZTCSt14basic_ifstreamIcSt11char_traitsIcEE0_Si RtlLookupFunctionEntry _ZGVNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr.__xi_a __imp_ungetwc _ZTINSt7__cxx118messagesIwEE _ZTCSt13basic_fstreamIcSt11char_traitsIcEE16_So _ZGVNSt10moneypunctIwLb0EE2idE __imp_fgetpos _ZTCSd0_Si _ZTISt8bad_cast _ZTISt9time_base _ZTSNSt7__cxx1115messages_bynameIwEE .refptr.__xi_z GetLastError __imp_ungetc _ZTINSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZTVSt10bad_typeid .refptr._ZTVSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE mingw_initltsdrot_force _head_lib64_libkernel32_a _ZGVNSt7collateIwE2idE _ZTISt9bad_alloc _ZTISt17__timepunct_cacheIwE .refptr._ZNSt8bad_castD1Ev _ZTI�	      St23__codecvt_abstract_baseIDsciE _ZNSt6locale5_Impl14_S_id_messagesE __imp_setvbuf __mingw_oldexcpt_handler _ZTISt23__codecvt_abstract_baseIwciE InitializeCriticalSection __imp_printf _ZTVSt14basic_ofstreamIcSt11char_traitsIcEE _ZTSNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE _ZTSNSt7__cxx1117moneypunct_bynameIwLb0EEE .refptr._ZSt7nothrow _ZTVSt14overflow_error _ZTSSt23__codecvt_abstract_baseIDiciE _tls_start _ZTISt17__timepunct_cacheIcE _ZTSSt7codecvtIwciE _ZTISt10money_base _ZTISt11range_error _ZTVN10__cxxabiv115__forced_unwindE _ZTSNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZTIN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE _ZNSt7__cxx1110moneypunctIwLb0EE2idE _ZTSN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE _ZNSt17moneypunct_bynameIwLb1EE4intlE __imp_GetCurrentProcessId _ZTISt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZNSt10__num_base11_S_atoms_inE _ZNSt6locale4noneE .refptr._ZNSt11__timepunctIwE2idE _ZT�	      VSt8messagesIcE __size_of_stack_reserve__ _ZTVNSt7__cxx1115numpunct_bynameIwEE .refptr._ZNSt10moneypunctIwLb1EE2idE _ZTINSt7__cxx1115numpunct_bynameIwEE _ZTSSt7codecvtIDiciE __getmainargs .refptr.__imp__acmdln _ZTVN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE __imp_putc _ZTSNSt7__cxx118numpunctIwEE _ZTSNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE __native_vcclrit_reason CreateEventA _ZNSt10moneypunctIwLb1EE4intlE _ZTISt16__numpunct_cacheIcE _ZTVNSt7__cxx1110moneypunctIwLb0EEE _ZTSNSt7__cxx1117moneypunct_bynameIcLb0EEE _ZTSSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZTVNSt7__cxx1115time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZTVNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEEE _ZTINSt7__cxx118numpunctIwEE _ZTSSt8numpunctIcE __imp___p__fmode _ZTCSt14basic_ofstreamIwSt11char_traitsIwEE0_St13basic_ostreamIwS1_E __imp_isspace _ZTVSt14collate_bynameIcE __imp__errno _ZNSt6locale5facet11_S_c_localeE __imp____lc_codepage�	      _func .refptr._ZN14__gnu_internal13buf_cout_syncE _ZNSt8ios_base3curE __imp_getchar _ZTINSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE ___lc_codepage_func _ZGVNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZTVSt13basic_filebufIcSt11char_traitsIcEE _ZTVSt14basic_iostreamIwSt11char_traitsIwEE __imp_CreateEventA __imp___p__acmdln __imp_exit _ZNSt7__cxx1117moneypunct_bynameIcLb1EE4intlE _ZTSSt25__codecvt_utf8_utf16_baseIwE _ZNSt6locale5_Impl19_S_facet_categoriesE _ZTISt7codecvtIcciE .refptr.mingw_app_type _ZTSN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE .refptr._ZNSt10moneypunctIcLb0EE2idE _ZTISt17moneypunct_bynameIcLb0EE .refptr._ZNSt7__cxx119money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt14basic_iostreamIwSt11char_traitsIwEE _ZTCSt14basic_ifstreamIwSt11char_traitsIwEE0_St13basic_istreamIwS1_E _ZSt4clog _ZTSNSt7__cxx1115messages_bynameIcEE DeleteCriticalSection SetLastError .refptr._ZN14__gnu_internal8buf_coutE .refptr.__imp___pioin�	      fo _ZTSNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE __imp__initterm _ZNSt10__num_base11_S_atoms_inE _ZNSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTSSt13basic_filebufIwSt11char_traitsIwEE __subsystem__ _ZTINSt8ios_base7failureB5cxx11E _ZTSSt8numpunctIwE _ZTISt20bad_array_new_length _ZTSSt14basic_ofstreamIwSt11char_traitsIwEE _ZTSSt15messages_bynameIcE _ZTVSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZSt5wclog __imp____mb_cur_max_func .refptr._ZNSt11__timepunctIcE2idE _ZTINSt7__cxx117collateIwEE __imp_fflush _ZTISt16__numpunct_cacheIwE _ZTCSt13basic_fstreamIwSt11char_traitsIwEE0_St14basic_iostreamIwS1_E _ZTTSt14basic_ifstreamIcSt11char_traitsIcEE _ZNSbIwSt11char_traitsIwESaIwEE4nposE .refptr._ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTIN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE __imp___C_specific_handler .refptr._ZTVNSt7__cxx119money_put�	      IcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEE .refptr._ZSt5wcout .refptr._ZN14__gnu_internal7buf_cinE __imp_GetCurrentProcess _ZTVSt23__codecvt_abstract_baseIDiciE __imp_MultiByteToWideChar _ZTISt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZGVNSt7__cxx118time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSbIwSt11char_traitsIwESaIwEE4_Rep20_S_empty_rep_storageE setlocale _ZTSNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .refptr._ZNSt7codecvtIcciE2idE _ZTSSt10ctype_base __imp_InitializeCriticalSection __lconv_init _filelengthi64 _ZTVNSt7__cxx118messagesIwEE .refptr._ZNSt6locale7_S_onceE ___crt_xi_start__ _ZNSt6locale10_S_classicE _ZNSt8ios_base5rightE _ZTSN9__gnu_cxx24__concurrence_wait_errorE _ZTVNSt7__cxx1115messages_bynameIcEE _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt23__codecvt_abstract_baseIcciE _ZNSs4_Rep20_S_empty_rep_storageE _ZTSSt17moneypunct_bynameIcLb0EE _lseeki64 .refptr._dowildcard __imp___doserrno _Z�	      TINSt7__cxx1117moneypunct_bynameIwLb0EEE _ZNSt8ios_base7unitbufE __imp__ultoa _ZTSSt18__moneypunct_cacheIcLb0EE _ZTSSt23__codecvt_abstract_baseIDsciE .refptr._ZTVSt10moneypunctIcLb1EE __imp__onexit __major_subsystem_version__ _ZTISt15messages_bynameIwE __bigtens_D2A _ZTSNSt7__cxx1110moneypunctIwLb1EEE _ZGVNSt8messagesIcE2idE _ZTVSt9basic_iosIwSt11char_traitsIwEE .refptr._ZNSt6locale13_S_categoriesE _ZTVSt23__codecvt_abstract_baseIcciE _ZTISt12ctype_bynameIwE _ZTSSt19__codecvt_utf8_baseIDsE _ZTVSt9bad_alloc _ZTVSt7codecvtIDsciE .refptr._ZNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZNSt5ctypeIcE2idE __imp_fopen .refptr._ZTVSt8numpunctIwE _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTSNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZTVNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZTVSt9type_info .refptr._ZNSt7collateIwE2idE _ZGVNSt8numpunctIcE2idE _ZTISt13runtime_error __mingw_winmain_hInstance __im�	      p_fclose __imp_ReleaseSemaphore _ZTISt17moneypunct_bynameIwLb0EE .refptr._ZNSt12out_of_rangeD1Ev _ZNSt8messagesIcE2idE _ZTIN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE MultiByteToWideChar ___crt_xt_end__ _ZTVSt20bad_array_new_length _ZTSSt20__codecvt_utf16_baseIDsE _ZNSt5ctypeIcE2idE TryEnterCriticalSection .refptr._ZTVSo RaiseException _ZTISt8ios_base .refptr._ZTVSt18__moneypunct_cacheIcLb1EE ___crt_xt_start__ _ZTSNSt3_V214error_categoryE .refptr._ZTVSi _ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt14collate_bynameIcE ___RUNTIME_PSEUDO_RELOC_LIST__ .refptr._ZTVSt23__codecvt_abstract_baseIwciE _ZTSSt10money_base .refptr.__mingw_oldexcpt_handler .refptr._ZTVSt10bad_typeid _ZGVNSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt13messages_base _ZTISt9type_info __imp_wcsftime _ZTSSt19__codecvt_utf8_baseIwE _ZTSSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSbIwSt11char_traitsIwESaIwEE4_Rep11_S_max_sizeE __imp___pioinfo __major_i�	      mage_version__ __section_alignment__ RtlAddFunctionTable .refptr._ZTVNSt7__cxx1110moneypunctIcLb1EEE _ZN14__gnu_internal13buf_cout_syncE _ZTINSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE .refptr._ZN10__cxxabiv120__unexpected_handlerE .refptr._ZSt4cout _ZTVSt19__codecvt_utf8_baseIDiE _ZTISt18__moneypunct_cacheIwLb0EE __imp_putwc __imp_GetSystemTimeAsFileTime _ZTVSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZTSNSt7__cxx1110moneypunctIcLb0EEE GetProcessAffinityMask _ZTISt7codecvtIDsciE _ZTSNSt7__cxx1115time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEE _ZTISt15messages_bynameIcE _ZTISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt10moneypunctIwLb1EE2idE .refptr.__native_startup_state _ZNSt10ctype_base5lowerE GetHandleInformation .refptr._ZNSt10moneypunctIcLb1EE2idE _ZTVSt17moneypunct_bynameIwLb0EE _ZTISt12codecvt_base ___crt_xl_start__ _ZNSt7codecvtIwciE2idE __DTOR_LIST__ _ZGVNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char�	      _traitsIcEEE2idE .refptr._ZNSt13runtime_errorD1Ev _ZSt5wclog _ZNSt10ctype_base5alphaE __imp_RtlCaptureContext _ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE GetTickCount __lib64_libmsvcrt_os_a_iname _ZTVSt17moneypunct_bynameIcLb1EE .refptr._ZTVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE _ZTSSt25__codecvt_utf8_utf16_baseIDiE _ZGVNSt11__timepunctIcE2idE __bss_start__ VirtualProtect _ZTVSt14basic_ofstreamIwSt11char_traitsIwEE mingw_initltsdyn_force .refptr._ZTVSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt19__iosfail_type_info _pthread_key_dest _ZNSt7__cxx1117moneypunct_bynameIwLb0EE4intlE _ZTVSt18__moneypunct_cacheIcLb0EE .refptr.__dyn_tls_init_callback .refptr._ZNSt7__cxx118messagesIwE2idE _ZTVNSt7__cxx1117moneypunct_bynameIcLb1EEE _ZTINSt6locale5facetE __minor_image_version__ _ZTVSt8numpunctIwE .refptr._ZTVSt15basic_streambufIcSt11char_traitsIcEE _ZTVNSt7__cxx1114collate_bynameIcEE .refptr._ZTVSt15basic_streambufIwSt11char_traitsIwEE .refptr�	      ._ZTVSt16__numpunct_cacheIwE mingw_initcharmax _ZTVSt12ctype_bynameIcE __imp_GetLastError _ZNSt10moneypunctIcLb1EE2idE _ZTVSt13basic_filebufIcSt11char_traitsIcEE UnhandledExceptionFilter _ZTSNSt7__cxx1117moneypunct_bynameIwLb1EEE _ZNSt8ios_base8showbaseE __imp_localeconv _ZNSt6locale8monetaryE _ZTVSt10moneypunctIwLb1EE ___crt_xp_end__ _ZNSt6locale2id11_S_refcountE __imp_VirtualProtect _ZNSt6locale5facet9_S_c_nameE _ZTCSt13basic_fstreamIwSt11char_traitsIwEE16_St13basic_ostreamIwS1_E _ZTVSt17__timepunct_cacheIwE _ZTSSt9basic_iosIcSt11char_traitsIcEE _ZGVNSt7__cxx1110moneypunctIcLb0EE2idE ___tls_start__ _ZGVNSt7__cxx119money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr._ZNSt20bad_array_new_lengthD1Ev _ZTSSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTSSt14basic_ifstreamIcSt11char_traitsIcEE _ZTVN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE _ZTISt14basic_ifstreamIwSt11char_traitsIwEE _ZTISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTTSt14basic_ifstr�	      eamIwSt11char_traitsIwEE .refptr.mingw_initltsdyn_force .refptr._ZTVSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZTVSt18__moneypunct_cacheIwLb0EE .refptr._ZNSt14overflow_errorD1Ev _ZNSt8ios_base9boolalphaE _ZTSNSt7__cxx1115numpunct_bynameIwEE _ZTSSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTSSt12ctype_bynameIwE __imp_strncmp _ZTSSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .refptr._ZTVSt15time_put_bynameIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE .refptr._ZNSt9bad_allocD1Ev _ZTISt10moneypunctIwLb0EE _ZTVNSt7__cxx1115messages_bynameIwEE _ZTSSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt8ios_base3decE __imp_TlsSetValue _ZNSt17__timepunct_cacheIwE12_S_timezonesE _ZTISt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE __mingw_pinit _MINGW_INSTALL_DEBUG_MATHERR _ZGVNSt7__cxx118messagesIwE2idE .refptr.__RUNTIME_PSEUDO_RELOC_LIST_END__ _tls_index __mingw_winmain_lpCmdLine __imp_getc _ZTSSt21__ctype_abstract_baseIcE _ZNSt�	      10moneypunctIcLb1EE4intlE _ZNSt10moneypunctIwLb0EE4intlE _ZTSSt13basic_istreamIwSt11char_traitsIwEE _ZNSt6locale7_S_onceE _ZNSt10ctype_base5blankE _ZTVNSt8ios_base7failureB5cxx11E .refptr._ZNSt8messagesIcE2idE _ZTVNSt7__cxx118numpunctIcEE .refptr._ZTVSt9bad_alloc __imp_memmove _ZNSt8ios_base3hexE .refptr.__tinytens_D2A _ZTISt21__ctype_abstract_baseIwE __IAT_start__ _ZTVSt12ctype_bynameIwE __imp_fputc _ZTSSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt19__codecvt_utf8_baseIDiE ___crt_xc_end__ __CTOR_LIST__ __setusermatherr _ZTSSt17moneypunct_bynameIwLb0EE _ZNSt7__cxx1110moneypunctIwLb1EE4intlE TlsSetValue __imp___iob_func __data_start__ _ZNSt7__cxx1117moneypunct_bynameIcLb0EE4intlE _ZNSt6locale17_S_twinned_facetsE _ZNSt8ios_base5fixedE _ZNSt8ios_base9basefieldE _ZNSt6locale9_S_globalE .refptr._ZTVSt13basic_filebufIwSt11char_traitsIwEE _initterm __imp_fwrite _ZTISt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZTVSt15time_get_bynameIwSt19istreambuf_iteratorIwSt11char_trait�	      sIwEEE _ZN14__gnu_internal12buf_cin_syncE _ZTVSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZNSt7__cxx117collateIcE2idE _ZTSSt17__timepunct_cacheIcE __imp_vfprintf _ZTCSt14basic_iostreamIwSt11char_traitsIwEE0_St13basic_istreamIwS1_E _ZTSNSt7__cxx118messagesIwEE _ZTVSt5ctypeIwE __imp_RtlUnwindEx _ZN14__gnu_internal8buf_wcinE __data_end__ WaitForMultipleObjects _ZTVSt14collate_bynameIwE _ZGVNSt7__cxx118numpunctIcE2idE _ZTSSt15basic_streambufIcSt11char_traitsIcEE _ZTSSt13runtime_error _ZTVSt13__ios_failure .refptr._ZTVSt16__numpunct_cacheIcE ___CTOR_LIST__ .refptr._ZNSt7codecvtIDiciE2idE __imp_ResumeThread _ZGVNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZN14__gnu_internal14buf_wcerr_syncE .refptr._ZTVSt14codecvt_bynameIcciE _ZGVNSt7__cxx118time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp_SetEvent _ZTTSt13basic_fstreamIcSt11char_traitsIcEE _ZTSSt16__numpunct_cacheIcE _ZNSt8ios_base3endE _ZTISt13basic_fstreamIcSt11char_traitsIcEE �	      _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt15basic_streambufIcSt11char_traitsIcEE _ZTSSt15underflow_error mingw_initltssuo_force __minor_os_version__ _ZNSt17moneypunct_bynameIcLb0EE4intlE __imp_TerminateProcess _ZTINSt7__cxx1115messages_bynameIcEE .refptr._ZN14__gnu_internal12buf_cin_syncE __imp__write __imp___initenv ___chkstk_ms .refptr._ZNSt15underflow_errorD1Ev _ZTISt25__codecvt_utf8_utf16_baseIDsE _ZTISt14codecvt_bynameIwciE .refptr._ZNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZTISt13basic_istreamIwSt11char_traitsIwEE _ZGVNSt7__cxx118messagesIcE2idE _ZTISt11__timepunctIwE _ZTSN10__cxxabiv119__foreign_exceptionE _ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZTVSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt5ctypeIcE10table_sizeE _ZTINSt7__cxx1117moneypunct_bynameIcLb0EEE _ZNSt7codecvtIDiciE2idE _ZTVSt8time_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE .refptr._ZTVNSt7__cxx119money_putIwSt1�	      9ostreambuf_iteratorIwSt11char_traitsIwEEEE __imp__fstat64 _ZTSSt8time_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE _ZTSSt9time_base _ZTVSt17__timepunct_cacheIcE .refptr._ZTVSt8bad_cast .refptr._ZTVSt11logic_error _ZTSN9__gnu_cxx24__concurrence_lock_errorE .refptr._ZNSt7__cxx119money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE .refptr._ZNSt7codecvtIwciE2idE _ZNSt6locale7numericE _ZSt5wcout _ZNSt10ctype_base6xdigitE _ZTSSt14overflow_error .refptr._ZTVNSt7__cxx117collateIwEE _ZTSSt14collate_bynameIwE _ZTINSt7__cxx118numpunctIcEE _ZNSt8ios_base3octE _ZGVNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZTISt14basic_ofstreamIcSt11char_traitsIcEE _ZTSNSt8ios_base7failureB5cxx11E _ZTTSt14basic_ofstreamIcSt11char_traitsIcEE .refptr._ZTVSt10moneypunctIwLb0EE _ZTVSt25__codecvt_utf8_utf16_baseIDsE __imp_realloc .refptr._ZTVSt13basic_istreamIwSt11char_traitsIwEE _ZTVSt5ctypeIcE .refptr.mingw_initltsdrot_force RtlCaptureContext _ZTSN9__gnu_cxx29__concurrence_broadcast_errorE _ZTVSt�	      20__codecvt_utf16_baseIDiE .refptr._ZTVNSt7__cxx1110moneypunctIwLb0EEE GetCurrentThreadId _ZTVNSt3_V214error_categoryE _ZTISt20__codecvt_utf16_baseIDsE _ZTSSt11logic_error _ZTVSt14codecvt_bynameIcciE _ZTVSt15messages_bynameIcE _ZTVSt13basic_ostreamIwSt11char_traitsIwEE __bss_end__ .refptr._ZTVSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE .refptr._ZTVSt5ctypeIcE _ZNSt7__cxx1110moneypunctIwLb0EE4intlE _ZTVSt21__ctype_abstract_baseIwE _ZNSt10moneypunctIcLb0EE4intlE _ZNSt7collateIwE2idE _ZNSt6locale7collateE __imp_fsetpos __imp_towupper _ZTSSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZNSt8ios_base4Init11_S_refcountE DuplicateHandle _ZNSbIwSt11char_traitsIwESaIwEE4_Rep11_S_terminalE _ZNSt9money_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZNSt7__cxx118numpunctIwE2idE _ZTVSt13basic_istreamIwSt11char_traitsIwEE .refptr._ZNSt11logic_errorD1Ev LeaveCriticalSection _ZTSSt14codecvt_bynameIwciE _ZTISt15numpunct_bynameIwE __ImageBase .refptr._ZNSt11range_errorD1Ev .refptr._ZT�	      VSt20bad_array_new_length .refptr._ZTVSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt8ios_base7goodbitE .refptr._ZTVSt9basic_iosIcSt11char_traitsIcEE _ZTVN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE __file_alignment__ _ZNSt8ios_base2inE .refptr._ZTVN9__gnu_cxx18stdio_sync_filebufIwSt11char_traitsIwEEE _ZTIN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE _ZTVSt11__timepunctIwE .refptr._ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZTISt9basic_iosIwSt11char_traitsIwEE _ZNSt7__cxx118messagesIwE2idE _ZTISt10moneypunctIcLb1EE __imp_strcmp _ZNSt7__cxx1110moneypunctIcLb0EE2idE _ZNSs4_Rep11_S_terminalE _ZTISt12out_of_range .refptr._ZN14__gnu_internal8buf_wcinE .refptr._ZTVSt18__moneypunct_cacheIwLb1EE .refptr._ZNSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE _ZGVNSt7num_putIwSt19ostreambuf_iteratorIwSt11char_traitsIwEEE2idE .refptr._ZTVSt9money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE _ZTVSt15underflow_error _ZTSSt15time_put_bynameIcSt19ostream�	      buf_iteratorIcSt11char_traitsIcEEE _ZTVSt10moneypunctIwLb0EE _ZSt5wcerr __imp_AddVectoredExceptionHandler _ZTISt14basic_ifstreamIcSt11char_traitsIcEE .refptr._ZTVSt13bad_exception _ZTVSt11__timepunctIcE .refptr._ZTVNSt7__cxx119money_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEEE .refptr._ZNSt8ios_base4Init20_S_synced_with_stdioE _ZTVNSt7__cxx1114collate_bynameIwEE _ZTSNSt7__cxx1115numpunct_bynameIcEE _ZGVNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt7__cxx1110moneypunctIcLb1EE4intlE _ZTSSt17__timepunct_cacheIwE .refptr._ZTVNSt7__cxx1110moneypunctIwLb1EEE _ZNSt8ios_base3appE _ZTSNSt6locale5facet6__shimE _ZTSSt8bad_cast __lib64_libkernel32_a_iname _ZNSt11__timepunctIcE2idE _ZTSSt10moneypunctIcLb1EE __imp_signal __dyn_tls_init_callback _ZTSSt14collate_bynameIcE .refptr._ZNSt7num_getIwSt19istreambuf_iteratorIwSt11char_traitsIwEEE2idE __imp_IsDBCSLeadByteEx GetSystemTimeAsFileTime __imp_UnhandledExceptionFilter .refptr._ZNSt8messagesIwE2idE _ZTVSt21__ctype_abstract_baseIcE _ZNS�	      t8ios_base7showposE __size_of_stack_commit__ _ZNSt7__cxx118numpunctIcE2idE RtlUnwindEx _ZTISt11__timepunctIcE _ZGVNSt10moneypunctIwLb1EE2idE __dll_characteristics__ _ZNSt10ctype_base5cntrlE .refptr.__native_startup_lock __imp__setjmp _ZTSN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE _ZTISt17moneypunct_bynameIwLb1EE __imp_memset _ZTSSt12ctype_bynameIcE __imp_ResetEvent _ZNSt6locale8messagesE _ZTSNSt8ios_base7failureE _ZNSt10ctype_base5punctE _ZTINSt7__cxx1117moneypunct_bynameIwLb1EEE _ZTSSt23__codecvt_abstract_baseIwciE _ZTISt23__codecvt_abstract_baseIDiciE _ZNSt8ios_base10floatfieldE _ZTISt8numpunctIcE _ZNSt8ios_base6skipwsE _ZTVSt23__codecvt_abstract_baseIwciE _ZTVSt23__codecvt_abstract_baseIDsciE _ZTSSt15messages_bynameIwE .refptr._ZNSt16invalid_argumentD1Ev _ZTISt15underflow_error _ZTSNSt6locale5facetE _ZTSSt10moneypunctIwLb1EE _ZGVNSt8messagesIwE2idE VirtualQuery _ZTISt14collate_bynameIwE _ZTVSt16__numpunct_cacheIcE __imp_strerror localeconv .refptr._ZNSt6locale17_S_twinned_facetsE _ZTVNSt7__cx�	      x1110moneypunctIcLb1EEE ze_of_stack_commit__ _ZNSt7__cxx118numpunctIcE2idE RtlUnwindEx _ZTISt11__timepunctIcE _ZGVNSt10moneypunctIwLb1EE2idE __dll_characteristics__ _ZNSt10ctype_base5cntrlE .refptr.__native_startup_lock __imp__setjmp _ZTSN9__gnu_cxx13stdio_filebufIwSt11char_traitsIwEEE _ZTISt17moneypunct_bynameIwLb1EE __imp_memset _ZTSSt12ctype_bynameIcE __imp_ResetEvent _ZNSt6locale8messagesE _ZTSNSt8ios_base7failureE _ZNSt10ctype_base5punctE _ZTINSt7__cxx1117moneypunct_bynameIwLb1EEE _ZTSSt23__codecvt_abstract_baseIwciE _ZTISt23__codecvt_abstract_baseIDiciE _ZNSt8ios_base10floatfieldE _ZTISt8numpunctIcE _ZNSt8ios_base6skipwsE _ZTVSt23__codecvt_abstract_baseIwciE _ZTVSt23__codecvt_abstract_baseIDsciE _ZTSSt15messages_bynameIwE .refptr._ZNSt16invalid_argumentD1Ev _ZTISt15underflow_error _ZTSNSt6locale5facetE _ZTSSt10moneypunctIwLb1EE _ZGVNSt8messagesIwE2idE VirtualQuery _ZTISt14collate_bynameIwE _ZTVSt16__numpunct_cacheIcE __imp_strerror localeconv .refptr._ZNSt6locale17_S_twinned_facetsE _ZTVNSt7__cx�	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              #                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              )                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              /                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              N                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              O                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              [                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ^                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              _                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              a                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              f                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              g                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              i                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              q                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              {                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              |                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              }                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
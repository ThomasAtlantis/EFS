	              � s��    s��    �     "�t��          I�t��                  8                                            0(r                    x      �      z       (r     �       (r     �      x             z                     8D���  p         ����@a�              a�           �      z      0(r     x        �    z             �     �      }       (r     z        �    }      �      � �   x      �              }      x      z {           z      �      �'r     �&r     � �    z      � �    }      }      x y           %r     �      z             � �           z {            � �    %�t��  � �       �  � �            � �     (r     � �              �     t�                  �$r     �'r      N}             �     t�    (              �$r             N}                  Ѓs�           �                      0(r     Ѓs��  �1R��         \�p     �$r     Y      Y�p            ��L��  �1R��              ڥ���  Y      ^�p     